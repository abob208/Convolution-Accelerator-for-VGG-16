`timescale 1ns / 1ns
module line_buffer ( clk, pixel_00, pixel_01, pixel_02, pixel_10, pixel_11, 
        pixel_12, pixel_20, pixel_21, pixel_22, in_pixel );
  output [7:0] pixel_00;
  output [7:0] pixel_01;
  output [7:0] pixel_02;
  output [7:0] pixel_10;
  output [7:0] pixel_11;
  output [7:0] pixel_12;
  output [7:0] pixel_20;
  output [7:0] pixel_21;
  output [7:0] pixel_22;
  input [7:0] in_pixel;
  input clk;
  wire   \row2_buffer[0][7] , \row2_buffer[0][6] , \row2_buffer[0][5] ,
         \row2_buffer[0][4] , \row2_buffer[0][3] , \row2_buffer[0][2] ,
         \row2_buffer[0][1] , \row2_buffer[0][0] , \row2_buffer[1][7] ,
         \row2_buffer[1][6] , \row2_buffer[1][5] , \row2_buffer[1][4] ,
         \row2_buffer[1][3] , \row2_buffer[1][2] , \row2_buffer[1][1] ,
         \row2_buffer[1][0] , \row2_buffer[2][7] , \row2_buffer[2][6] ,
         \row2_buffer[2][5] , \row2_buffer[2][4] , \row2_buffer[2][3] ,
         \row2_buffer[2][2] , \row2_buffer[2][1] , \row2_buffer[2][0] ,
         \row2_buffer[3][7] , \row2_buffer[3][6] , \row2_buffer[3][5] ,
         \row2_buffer[3][4] , \row2_buffer[3][3] , \row2_buffer[3][2] ,
         \row2_buffer[3][1] , \row2_buffer[3][0] , \row2_buffer[4][7] ,
         \row2_buffer[4][6] , \row2_buffer[4][5] , \row2_buffer[4][4] ,
         \row2_buffer[4][3] , \row2_buffer[4][2] , \row2_buffer[4][1] ,
         \row2_buffer[4][0] , \row2_buffer[5][7] , \row2_buffer[5][6] ,
         \row2_buffer[5][5] , \row2_buffer[5][4] , \row2_buffer[5][3] ,
         \row2_buffer[5][2] , \row2_buffer[5][1] , \row2_buffer[5][0] ,
         \row2_buffer[6][7] , \row2_buffer[6][6] , \row2_buffer[6][5] ,
         \row2_buffer[6][4] , \row2_buffer[6][3] , \row2_buffer[6][2] ,
         \row2_buffer[6][1] , \row2_buffer[6][0] , \row2_buffer[7][7] ,
         \row2_buffer[7][6] , \row2_buffer[7][5] , \row2_buffer[7][4] ,
         \row2_buffer[7][3] , \row2_buffer[7][2] , \row2_buffer[7][1] ,
         \row2_buffer[7][0] , \row2_buffer[8][7] , \row2_buffer[8][6] ,
         \row2_buffer[8][5] , \row2_buffer[8][4] , \row2_buffer[8][3] ,
         \row2_buffer[8][2] , \row2_buffer[8][1] , \row2_buffer[8][0] ,
         \row2_buffer[9][7] , \row2_buffer[9][6] , \row2_buffer[9][5] ,
         \row2_buffer[9][4] , \row2_buffer[9][3] , \row2_buffer[9][2] ,
         \row2_buffer[9][1] , \row2_buffer[9][0] , \row2_buffer[10][7] ,
         \row2_buffer[10][6] , \row2_buffer[10][5] , \row2_buffer[10][4] ,
         \row2_buffer[10][3] , \row2_buffer[10][2] , \row2_buffer[10][1] ,
         \row2_buffer[10][0] , \row2_buffer[11][7] , \row2_buffer[11][6] ,
         \row2_buffer[11][5] , \row2_buffer[11][4] , \row2_buffer[11][3] ,
         \row2_buffer[11][2] , \row2_buffer[11][1] , \row2_buffer[11][0] ,
         \row2_buffer[12][7] , \row2_buffer[12][6] , \row2_buffer[12][5] ,
         \row2_buffer[12][4] , \row2_buffer[12][3] , \row2_buffer[12][2] ,
         \row2_buffer[12][1] , \row2_buffer[12][0] , \row2_buffer[13][7] ,
         \row2_buffer[13][6] , \row2_buffer[13][5] , \row2_buffer[13][4] ,
         \row2_buffer[13][3] , \row2_buffer[13][2] , \row2_buffer[13][1] ,
         \row2_buffer[13][0] , \row2_buffer[14][7] , \row2_buffer[14][6] ,
         \row2_buffer[14][5] , \row2_buffer[14][4] , \row2_buffer[14][3] ,
         \row2_buffer[14][2] , \row2_buffer[14][1] , \row2_buffer[14][0] ,
         \row2_buffer[15][7] , \row2_buffer[15][6] , \row2_buffer[15][5] ,
         \row2_buffer[15][4] , \row2_buffer[15][3] , \row2_buffer[15][2] ,
         \row2_buffer[15][1] , \row2_buffer[15][0] , \row2_buffer[16][7] ,
         \row2_buffer[16][6] , \row2_buffer[16][5] , \row2_buffer[16][4] ,
         \row2_buffer[16][3] , \row2_buffer[16][2] , \row2_buffer[16][1] ,
         \row2_buffer[16][0] , \row2_buffer[17][7] , \row2_buffer[17][6] ,
         \row2_buffer[17][5] , \row2_buffer[17][4] , \row2_buffer[17][3] ,
         \row2_buffer[17][2] , \row2_buffer[17][1] , \row2_buffer[17][0] ,
         \row2_buffer[18][7] , \row2_buffer[18][6] , \row2_buffer[18][5] ,
         \row2_buffer[18][4] , \row2_buffer[18][3] , \row2_buffer[18][2] ,
         \row2_buffer[18][1] , \row2_buffer[18][0] , \row2_buffer[19][7] ,
         \row2_buffer[19][6] , \row2_buffer[19][5] , \row2_buffer[19][4] ,
         \row2_buffer[19][3] , \row2_buffer[19][2] , \row2_buffer[19][1] ,
         \row2_buffer[19][0] , \row2_buffer[20][7] , \row2_buffer[20][6] ,
         \row2_buffer[20][5] , \row2_buffer[20][4] , \row2_buffer[20][3] ,
         \row2_buffer[20][2] , \row2_buffer[20][1] , \row2_buffer[20][0] ,
         \row2_buffer[21][7] , \row2_buffer[21][6] , \row2_buffer[21][5] ,
         \row2_buffer[21][4] , \row2_buffer[21][3] , \row2_buffer[21][2] ,
         \row2_buffer[21][1] , \row2_buffer[21][0] , \row2_buffer[22][7] ,
         \row2_buffer[22][6] , \row2_buffer[22][5] , \row2_buffer[22][4] ,
         \row2_buffer[22][3] , \row2_buffer[22][2] , \row2_buffer[22][1] ,
         \row2_buffer[22][0] , \row2_buffer[23][7] , \row2_buffer[23][6] ,
         \row2_buffer[23][5] , \row2_buffer[23][4] , \row2_buffer[23][3] ,
         \row2_buffer[23][2] , \row2_buffer[23][1] , \row2_buffer[23][0] ,
         \row2_buffer[24][7] , \row2_buffer[24][6] , \row2_buffer[24][5] ,
         \row2_buffer[24][4] , \row2_buffer[24][3] , \row2_buffer[24][2] ,
         \row2_buffer[24][1] , \row2_buffer[24][0] , \row2_buffer[25][7] ,
         \row2_buffer[25][6] , \row2_buffer[25][5] , \row2_buffer[25][4] ,
         \row2_buffer[25][3] , \row2_buffer[25][2] , \row2_buffer[25][1] ,
         \row2_buffer[25][0] , \row2_buffer[26][7] , \row2_buffer[26][6] ,
         \row2_buffer[26][5] , \row2_buffer[26][4] , \row2_buffer[26][3] ,
         \row2_buffer[26][2] , \row2_buffer[26][1] , \row2_buffer[26][0] ,
         \row2_buffer[27][7] , \row2_buffer[27][6] , \row2_buffer[27][5] ,
         \row2_buffer[27][4] , \row2_buffer[27][3] , \row2_buffer[27][2] ,
         \row2_buffer[27][1] , \row2_buffer[27][0] , \row2_buffer[28][7] ,
         \row2_buffer[28][6] , \row2_buffer[28][5] , \row2_buffer[28][4] ,
         \row2_buffer[28][3] , \row2_buffer[28][2] , \row2_buffer[28][1] ,
         \row2_buffer[28][0] , \row2_buffer[29][7] , \row2_buffer[29][6] ,
         \row2_buffer[29][5] , \row2_buffer[29][4] , \row2_buffer[29][3] ,
         \row2_buffer[29][2] , \row2_buffer[29][1] , \row2_buffer[29][0] ,
         \row2_buffer[30][7] , \row2_buffer[30][6] , \row2_buffer[30][5] ,
         \row2_buffer[30][4] , \row2_buffer[30][3] , \row2_buffer[30][2] ,
         \row2_buffer[30][1] , \row2_buffer[30][0] , \row2_buffer[31][7] ,
         \row2_buffer[31][6] , \row2_buffer[31][5] , \row2_buffer[31][4] ,
         \row2_buffer[31][3] , \row2_buffer[31][2] , \row2_buffer[31][1] ,
         \row2_buffer[31][0] , \row2_buffer[32][7] , \row2_buffer[32][6] ,
         \row2_buffer[32][5] , \row2_buffer[32][4] , \row2_buffer[32][3] ,
         \row2_buffer[32][2] , \row2_buffer[32][1] , \row2_buffer[32][0] ,
         \row2_buffer[33][7] , \row2_buffer[33][6] , \row2_buffer[33][5] ,
         \row2_buffer[33][4] , \row2_buffer[33][3] , \row2_buffer[33][2] ,
         \row2_buffer[33][1] , \row2_buffer[33][0] , \row2_buffer[34][7] ,
         \row2_buffer[34][6] , \row2_buffer[34][5] , \row2_buffer[34][4] ,
         \row2_buffer[34][3] , \row2_buffer[34][2] , \row2_buffer[34][1] ,
         \row2_buffer[34][0] , \row2_buffer[35][7] , \row2_buffer[35][6] ,
         \row2_buffer[35][5] , \row2_buffer[35][4] , \row2_buffer[35][3] ,
         \row2_buffer[35][2] , \row2_buffer[35][1] , \row2_buffer[35][0] ,
         \row2_buffer[36][7] , \row2_buffer[36][6] , \row2_buffer[36][5] ,
         \row2_buffer[36][4] , \row2_buffer[36][3] , \row2_buffer[36][2] ,
         \row2_buffer[36][1] , \row2_buffer[36][0] , \row2_buffer[37][7] ,
         \row2_buffer[37][6] , \row2_buffer[37][5] , \row2_buffer[37][4] ,
         \row2_buffer[37][3] , \row2_buffer[37][2] , \row2_buffer[37][1] ,
         \row2_buffer[37][0] , \row2_buffer[38][7] , \row2_buffer[38][6] ,
         \row2_buffer[38][5] , \row2_buffer[38][4] , \row2_buffer[38][3] ,
         \row2_buffer[38][2] , \row2_buffer[38][1] , \row2_buffer[38][0] ,
         \row2_buffer[39][7] , \row2_buffer[39][6] , \row2_buffer[39][5] ,
         \row2_buffer[39][4] , \row2_buffer[39][3] , \row2_buffer[39][2] ,
         \row2_buffer[39][1] , \row2_buffer[39][0] , \row2_buffer[40][7] ,
         \row2_buffer[40][6] , \row2_buffer[40][5] , \row2_buffer[40][4] ,
         \row2_buffer[40][3] , \row2_buffer[40][2] , \row2_buffer[40][1] ,
         \row2_buffer[40][0] , \row2_buffer[41][7] , \row2_buffer[41][6] ,
         \row2_buffer[41][5] , \row2_buffer[41][4] , \row2_buffer[41][3] ,
         \row2_buffer[41][2] , \row2_buffer[41][1] , \row2_buffer[41][0] ,
         \row2_buffer[42][7] , \row2_buffer[42][6] , \row2_buffer[42][5] ,
         \row2_buffer[42][4] , \row2_buffer[42][3] , \row2_buffer[42][2] ,
         \row2_buffer[42][1] , \row2_buffer[42][0] , \row2_buffer[43][7] ,
         \row2_buffer[43][6] , \row2_buffer[43][5] , \row2_buffer[43][4] ,
         \row2_buffer[43][3] , \row2_buffer[43][2] , \row2_buffer[43][1] ,
         \row2_buffer[43][0] , \row2_buffer[44][7] , \row2_buffer[44][6] ,
         \row2_buffer[44][5] , \row2_buffer[44][4] , \row2_buffer[44][3] ,
         \row2_buffer[44][2] , \row2_buffer[44][1] , \row2_buffer[44][0] ,
         \row2_buffer[45][7] , \row2_buffer[45][6] , \row2_buffer[45][5] ,
         \row2_buffer[45][4] , \row2_buffer[45][3] , \row2_buffer[45][2] ,
         \row2_buffer[45][1] , \row2_buffer[45][0] , \row2_buffer[46][7] ,
         \row2_buffer[46][6] , \row2_buffer[46][5] , \row2_buffer[46][4] ,
         \row2_buffer[46][3] , \row2_buffer[46][2] , \row2_buffer[46][1] ,
         \row2_buffer[46][0] , \row2_buffer[47][7] , \row2_buffer[47][6] ,
         \row2_buffer[47][5] , \row2_buffer[47][4] , \row2_buffer[47][3] ,
         \row2_buffer[47][2] , \row2_buffer[47][1] , \row2_buffer[47][0] ,
         \row2_buffer[48][7] , \row2_buffer[48][6] , \row2_buffer[48][5] ,
         \row2_buffer[48][4] , \row2_buffer[48][3] , \row2_buffer[48][2] ,
         \row2_buffer[48][1] , \row2_buffer[48][0] , \row2_buffer[49][7] ,
         \row2_buffer[49][6] , \row2_buffer[49][5] , \row2_buffer[49][4] ,
         \row2_buffer[49][3] , \row2_buffer[49][2] , \row2_buffer[49][1] ,
         \row2_buffer[49][0] , \row2_buffer[50][7] , \row2_buffer[50][6] ,
         \row2_buffer[50][5] , \row2_buffer[50][4] , \row2_buffer[50][3] ,
         \row2_buffer[50][2] , \row2_buffer[50][1] , \row2_buffer[50][0] ,
         \row2_buffer[51][7] , \row2_buffer[51][6] , \row2_buffer[51][5] ,
         \row2_buffer[51][4] , \row2_buffer[51][3] , \row2_buffer[51][2] ,
         \row2_buffer[51][1] , \row2_buffer[51][0] , \row2_buffer[52][7] ,
         \row2_buffer[52][6] , \row2_buffer[52][5] , \row2_buffer[52][4] ,
         \row2_buffer[52][3] , \row2_buffer[52][2] , \row2_buffer[52][1] ,
         \row2_buffer[52][0] , \row2_buffer[53][7] , \row2_buffer[53][6] ,
         \row2_buffer[53][5] , \row2_buffer[53][4] , \row2_buffer[53][3] ,
         \row2_buffer[53][2] , \row2_buffer[53][1] , \row2_buffer[53][0] ,
         \row2_buffer[54][7] , \row2_buffer[54][6] , \row2_buffer[54][5] ,
         \row2_buffer[54][4] , \row2_buffer[54][3] , \row2_buffer[54][2] ,
         \row2_buffer[54][1] , \row2_buffer[54][0] , \row2_buffer[55][7] ,
         \row2_buffer[55][6] , \row2_buffer[55][5] , \row2_buffer[55][4] ,
         \row2_buffer[55][3] , \row2_buffer[55][2] , \row2_buffer[55][1] ,
         \row2_buffer[55][0] , \row2_buffer[56][7] , \row2_buffer[56][6] ,
         \row2_buffer[56][5] , \row2_buffer[56][4] , \row2_buffer[56][3] ,
         \row2_buffer[56][2] , \row2_buffer[56][1] , \row2_buffer[56][0] ,
         \row2_buffer[57][7] , \row2_buffer[57][6] , \row2_buffer[57][5] ,
         \row2_buffer[57][4] , \row2_buffer[57][3] , \row2_buffer[57][2] ,
         \row2_buffer[57][1] , \row2_buffer[57][0] , \row2_buffer[58][7] ,
         \row2_buffer[58][6] , \row2_buffer[58][5] , \row2_buffer[58][4] ,
         \row2_buffer[58][3] , \row2_buffer[58][2] , \row2_buffer[58][1] ,
         \row2_buffer[58][0] , \row2_buffer[59][7] , \row2_buffer[59][6] ,
         \row2_buffer[59][5] , \row2_buffer[59][4] , \row2_buffer[59][3] ,
         \row2_buffer[59][2] , \row2_buffer[59][1] , \row2_buffer[59][0] ,
         \row2_buffer[60][7] , \row2_buffer[60][6] , \row2_buffer[60][5] ,
         \row2_buffer[60][4] , \row2_buffer[60][3] , \row2_buffer[60][2] ,
         \row2_buffer[60][1] , \row2_buffer[60][0] , \row2_buffer[61][7] ,
         \row2_buffer[61][6] , \row2_buffer[61][5] , \row2_buffer[61][4] ,
         \row2_buffer[61][3] , \row2_buffer[61][2] , \row2_buffer[61][1] ,
         \row2_buffer[61][0] , \row2_buffer[62][7] , \row2_buffer[62][6] ,
         \row2_buffer[62][5] , \row2_buffer[62][4] , \row2_buffer[62][3] ,
         \row2_buffer[62][2] , \row2_buffer[62][1] , \row2_buffer[62][0] ,
         \row2_buffer[63][7] , \row2_buffer[63][6] , \row2_buffer[63][5] ,
         \row2_buffer[63][4] , \row2_buffer[63][3] , \row2_buffer[63][2] ,
         \row2_buffer[63][1] , \row2_buffer[63][0] , \row2_buffer[64][7] ,
         \row2_buffer[64][6] , \row2_buffer[64][5] , \row2_buffer[64][4] ,
         \row2_buffer[64][3] , \row2_buffer[64][2] , \row2_buffer[64][1] ,
         \row2_buffer[64][0] , \row2_buffer[65][7] , \row2_buffer[65][6] ,
         \row2_buffer[65][5] , \row2_buffer[65][4] , \row2_buffer[65][3] ,
         \row2_buffer[65][2] , \row2_buffer[65][1] , \row2_buffer[65][0] ,
         \row2_buffer[66][7] , \row2_buffer[66][6] , \row2_buffer[66][5] ,
         \row2_buffer[66][4] , \row2_buffer[66][3] , \row2_buffer[66][2] ,
         \row2_buffer[66][1] , \row2_buffer[66][0] , \row2_buffer[67][7] ,
         \row2_buffer[67][6] , \row2_buffer[67][5] , \row2_buffer[67][4] ,
         \row2_buffer[67][3] , \row2_buffer[67][2] , \row2_buffer[67][1] ,
         \row2_buffer[67][0] , \row2_buffer[68][7] , \row2_buffer[68][6] ,
         \row2_buffer[68][5] , \row2_buffer[68][4] , \row2_buffer[68][3] ,
         \row2_buffer[68][2] , \row2_buffer[68][1] , \row2_buffer[68][0] ,
         \row2_buffer[69][7] , \row2_buffer[69][6] , \row2_buffer[69][5] ,
         \row2_buffer[69][4] , \row2_buffer[69][3] , \row2_buffer[69][2] ,
         \row2_buffer[69][1] , \row2_buffer[69][0] , \row2_buffer[70][7] ,
         \row2_buffer[70][6] , \row2_buffer[70][5] , \row2_buffer[70][4] ,
         \row2_buffer[70][3] , \row2_buffer[70][2] , \row2_buffer[70][1] ,
         \row2_buffer[70][0] , \row2_buffer[71][7] , \row2_buffer[71][6] ,
         \row2_buffer[71][5] , \row2_buffer[71][4] , \row2_buffer[71][3] ,
         \row2_buffer[71][2] , \row2_buffer[71][1] , \row2_buffer[71][0] ,
         \row2_buffer[72][7] , \row2_buffer[72][6] , \row2_buffer[72][5] ,
         \row2_buffer[72][4] , \row2_buffer[72][3] , \row2_buffer[72][2] ,
         \row2_buffer[72][1] , \row2_buffer[72][0] , \row2_buffer[73][7] ,
         \row2_buffer[73][6] , \row2_buffer[73][5] , \row2_buffer[73][4] ,
         \row2_buffer[73][3] , \row2_buffer[73][2] , \row2_buffer[73][1] ,
         \row2_buffer[73][0] , \row2_buffer[74][7] , \row2_buffer[74][6] ,
         \row2_buffer[74][5] , \row2_buffer[74][4] , \row2_buffer[74][3] ,
         \row2_buffer[74][2] , \row2_buffer[74][1] , \row2_buffer[74][0] ,
         \row2_buffer[75][7] , \row2_buffer[75][6] , \row2_buffer[75][5] ,
         \row2_buffer[75][4] , \row2_buffer[75][3] , \row2_buffer[75][2] ,
         \row2_buffer[75][1] , \row2_buffer[75][0] , \row2_buffer[76][7] ,
         \row2_buffer[76][6] , \row2_buffer[76][5] , \row2_buffer[76][4] ,
         \row2_buffer[76][3] , \row2_buffer[76][2] , \row2_buffer[76][1] ,
         \row2_buffer[76][0] , \row2_buffer[77][7] , \row2_buffer[77][6] ,
         \row2_buffer[77][5] , \row2_buffer[77][4] , \row2_buffer[77][3] ,
         \row2_buffer[77][2] , \row2_buffer[77][1] , \row2_buffer[77][0] ,
         \row2_buffer[78][7] , \row2_buffer[78][6] , \row2_buffer[78][5] ,
         \row2_buffer[78][4] , \row2_buffer[78][3] , \row2_buffer[78][2] ,
         \row2_buffer[78][1] , \row2_buffer[78][0] , \row2_buffer[79][7] ,
         \row2_buffer[79][6] , \row2_buffer[79][5] , \row2_buffer[79][4] ,
         \row2_buffer[79][3] , \row2_buffer[79][2] , \row2_buffer[79][1] ,
         \row2_buffer[79][0] , \row2_buffer[80][7] , \row2_buffer[80][6] ,
         \row2_buffer[80][5] , \row2_buffer[80][4] , \row2_buffer[80][3] ,
         \row2_buffer[80][2] , \row2_buffer[80][1] , \row2_buffer[80][0] ,
         \row2_buffer[81][7] , \row2_buffer[81][6] , \row2_buffer[81][5] ,
         \row2_buffer[81][4] , \row2_buffer[81][3] , \row2_buffer[81][2] ,
         \row2_buffer[81][1] , \row2_buffer[81][0] , \row2_buffer[82][7] ,
         \row2_buffer[82][6] , \row2_buffer[82][5] , \row2_buffer[82][4] ,
         \row2_buffer[82][3] , \row2_buffer[82][2] , \row2_buffer[82][1] ,
         \row2_buffer[82][0] , \row2_buffer[83][7] , \row2_buffer[83][6] ,
         \row2_buffer[83][5] , \row2_buffer[83][4] , \row2_buffer[83][3] ,
         \row2_buffer[83][2] , \row2_buffer[83][1] , \row2_buffer[83][0] ,
         \row2_buffer[84][7] , \row2_buffer[84][6] , \row2_buffer[84][5] ,
         \row2_buffer[84][4] , \row2_buffer[84][3] , \row2_buffer[84][2] ,
         \row2_buffer[84][1] , \row2_buffer[84][0] , \row2_buffer[85][7] ,
         \row2_buffer[85][6] , \row2_buffer[85][5] , \row2_buffer[85][4] ,
         \row2_buffer[85][3] , \row2_buffer[85][2] , \row2_buffer[85][1] ,
         \row2_buffer[85][0] , \row2_buffer[86][7] , \row2_buffer[86][6] ,
         \row2_buffer[86][5] , \row2_buffer[86][4] , \row2_buffer[86][3] ,
         \row2_buffer[86][2] , \row2_buffer[86][1] , \row2_buffer[86][0] ,
         \row2_buffer[87][7] , \row2_buffer[87][6] , \row2_buffer[87][5] ,
         \row2_buffer[87][4] , \row2_buffer[87][3] , \row2_buffer[87][2] ,
         \row2_buffer[87][1] , \row2_buffer[87][0] , \row2_buffer[88][7] ,
         \row2_buffer[88][6] , \row2_buffer[88][5] , \row2_buffer[88][4] ,
         \row2_buffer[88][3] , \row2_buffer[88][2] , \row2_buffer[88][1] ,
         \row2_buffer[88][0] , \row2_buffer[89][7] , \row2_buffer[89][6] ,
         \row2_buffer[89][5] , \row2_buffer[89][4] , \row2_buffer[89][3] ,
         \row2_buffer[89][2] , \row2_buffer[89][1] , \row2_buffer[89][0] ,
         \row2_buffer[90][7] , \row2_buffer[90][6] , \row2_buffer[90][5] ,
         \row2_buffer[90][4] , \row2_buffer[90][3] , \row2_buffer[90][2] ,
         \row2_buffer[90][1] , \row2_buffer[90][0] , \row2_buffer[91][7] ,
         \row2_buffer[91][6] , \row2_buffer[91][5] , \row2_buffer[91][4] ,
         \row2_buffer[91][3] , \row2_buffer[91][2] , \row2_buffer[91][1] ,
         \row2_buffer[91][0] , \row2_buffer[92][7] , \row2_buffer[92][6] ,
         \row2_buffer[92][5] , \row2_buffer[92][4] , \row2_buffer[92][3] ,
         \row2_buffer[92][2] , \row2_buffer[92][1] , \row2_buffer[92][0] ,
         \row2_buffer[93][7] , \row2_buffer[93][6] , \row2_buffer[93][5] ,
         \row2_buffer[93][4] , \row2_buffer[93][3] , \row2_buffer[93][2] ,
         \row2_buffer[93][1] , \row2_buffer[93][0] , \row2_buffer[94][7] ,
         \row2_buffer[94][6] , \row2_buffer[94][5] , \row2_buffer[94][4] ,
         \row2_buffer[94][3] , \row2_buffer[94][2] , \row2_buffer[94][1] ,
         \row2_buffer[94][0] , \row2_buffer[95][7] , \row2_buffer[95][6] ,
         \row2_buffer[95][5] , \row2_buffer[95][4] , \row2_buffer[95][3] ,
         \row2_buffer[95][2] , \row2_buffer[95][1] , \row2_buffer[95][0] ,
         \row2_buffer[96][7] , \row2_buffer[96][6] , \row2_buffer[96][5] ,
         \row2_buffer[96][4] , \row2_buffer[96][3] , \row2_buffer[96][2] ,
         \row2_buffer[96][1] , \row2_buffer[96][0] , \row2_buffer[97][7] ,
         \row2_buffer[97][6] , \row2_buffer[97][5] , \row2_buffer[97][4] ,
         \row2_buffer[97][3] , \row2_buffer[97][2] , \row2_buffer[97][1] ,
         \row2_buffer[97][0] , \row2_buffer[98][7] , \row2_buffer[98][6] ,
         \row2_buffer[98][5] , \row2_buffer[98][4] , \row2_buffer[98][3] ,
         \row2_buffer[98][2] , \row2_buffer[98][1] , \row2_buffer[98][0] ,
         \row2_buffer[99][7] , \row2_buffer[99][6] , \row2_buffer[99][5] ,
         \row2_buffer[99][4] , \row2_buffer[99][3] , \row2_buffer[99][2] ,
         \row2_buffer[99][1] , \row2_buffer[99][0] , \row2_buffer[100][7] ,
         \row2_buffer[100][6] , \row2_buffer[100][5] , \row2_buffer[100][4] ,
         \row2_buffer[100][3] , \row2_buffer[100][2] , \row2_buffer[100][1] ,
         \row2_buffer[100][0] , \row2_buffer[101][7] , \row2_buffer[101][6] ,
         \row2_buffer[101][5] , \row2_buffer[101][4] , \row2_buffer[101][3] ,
         \row2_buffer[101][2] , \row2_buffer[101][1] , \row2_buffer[101][0] ,
         \row2_buffer[102][7] , \row2_buffer[102][6] , \row2_buffer[102][5] ,
         \row2_buffer[102][4] , \row2_buffer[102][3] , \row2_buffer[102][2] ,
         \row2_buffer[102][1] , \row2_buffer[102][0] , \row2_buffer[103][7] ,
         \row2_buffer[103][6] , \row2_buffer[103][5] , \row2_buffer[103][4] ,
         \row2_buffer[103][3] , \row2_buffer[103][2] , \row2_buffer[103][1] ,
         \row2_buffer[103][0] , \row2_buffer[104][7] , \row2_buffer[104][6] ,
         \row2_buffer[104][5] , \row2_buffer[104][4] , \row2_buffer[104][3] ,
         \row2_buffer[104][2] , \row2_buffer[104][1] , \row2_buffer[104][0] ,
         \row2_buffer[105][7] , \row2_buffer[105][6] , \row2_buffer[105][5] ,
         \row2_buffer[105][4] , \row2_buffer[105][3] , \row2_buffer[105][2] ,
         \row2_buffer[105][1] , \row2_buffer[105][0] , \row2_buffer[106][7] ,
         \row2_buffer[106][6] , \row2_buffer[106][5] , \row2_buffer[106][4] ,
         \row2_buffer[106][3] , \row2_buffer[106][2] , \row2_buffer[106][1] ,
         \row2_buffer[106][0] , \row2_buffer[107][7] , \row2_buffer[107][6] ,
         \row2_buffer[107][5] , \row2_buffer[107][4] , \row2_buffer[107][3] ,
         \row2_buffer[107][2] , \row2_buffer[107][1] , \row2_buffer[107][0] ,
         \row2_buffer[108][7] , \row2_buffer[108][6] , \row2_buffer[108][5] ,
         \row2_buffer[108][4] , \row2_buffer[108][3] , \row2_buffer[108][2] ,
         \row2_buffer[108][1] , \row2_buffer[108][0] , \row2_buffer[109][7] ,
         \row2_buffer[109][6] , \row2_buffer[109][5] , \row2_buffer[109][4] ,
         \row2_buffer[109][3] , \row2_buffer[109][2] , \row2_buffer[109][1] ,
         \row2_buffer[109][0] , \row2_buffer[110][7] , \row2_buffer[110][6] ,
         \row2_buffer[110][5] , \row2_buffer[110][4] , \row2_buffer[110][3] ,
         \row2_buffer[110][2] , \row2_buffer[110][1] , \row2_buffer[110][0] ,
         \row2_buffer[111][7] , \row2_buffer[111][6] , \row2_buffer[111][5] ,
         \row2_buffer[111][4] , \row2_buffer[111][3] , \row2_buffer[111][2] ,
         \row2_buffer[111][1] , \row2_buffer[111][0] , \row2_buffer[112][7] ,
         \row2_buffer[112][6] , \row2_buffer[112][5] , \row2_buffer[112][4] ,
         \row2_buffer[112][3] , \row2_buffer[112][2] , \row2_buffer[112][1] ,
         \row2_buffer[112][0] , \row2_buffer[113][7] , \row2_buffer[113][6] ,
         \row2_buffer[113][5] , \row2_buffer[113][4] , \row2_buffer[113][3] ,
         \row2_buffer[113][2] , \row2_buffer[113][1] , \row2_buffer[113][0] ,
         \row2_buffer[114][7] , \row2_buffer[114][6] , \row2_buffer[114][5] ,
         \row2_buffer[114][4] , \row2_buffer[114][3] , \row2_buffer[114][2] ,
         \row2_buffer[114][1] , \row2_buffer[114][0] , \row2_buffer[115][7] ,
         \row2_buffer[115][6] , \row2_buffer[115][5] , \row2_buffer[115][4] ,
         \row2_buffer[115][3] , \row2_buffer[115][2] , \row2_buffer[115][1] ,
         \row2_buffer[115][0] , \row2_buffer[116][7] , \row2_buffer[116][6] ,
         \row2_buffer[116][5] , \row2_buffer[116][4] , \row2_buffer[116][3] ,
         \row2_buffer[116][2] , \row2_buffer[116][1] , \row2_buffer[116][0] ,
         \row2_buffer[117][7] , \row2_buffer[117][6] , \row2_buffer[117][5] ,
         \row2_buffer[117][4] , \row2_buffer[117][3] , \row2_buffer[117][2] ,
         \row2_buffer[117][1] , \row2_buffer[117][0] , \row2_buffer[118][7] ,
         \row2_buffer[118][6] , \row2_buffer[118][5] , \row2_buffer[118][4] ,
         \row2_buffer[118][3] , \row2_buffer[118][2] , \row2_buffer[118][1] ,
         \row2_buffer[118][0] , \row2_buffer[119][7] , \row2_buffer[119][6] ,
         \row2_buffer[119][5] , \row2_buffer[119][4] , \row2_buffer[119][3] ,
         \row2_buffer[119][2] , \row2_buffer[119][1] , \row2_buffer[119][0] ,
         \row2_buffer[120][7] , \row2_buffer[120][6] , \row2_buffer[120][5] ,
         \row2_buffer[120][4] , \row2_buffer[120][3] , \row2_buffer[120][2] ,
         \row2_buffer[120][1] , \row2_buffer[120][0] , \row2_buffer[121][7] ,
         \row2_buffer[121][6] , \row2_buffer[121][5] , \row2_buffer[121][4] ,
         \row2_buffer[121][3] , \row2_buffer[121][2] , \row2_buffer[121][1] ,
         \row2_buffer[121][0] , \row2_buffer[122][7] , \row2_buffer[122][6] ,
         \row2_buffer[122][5] , \row2_buffer[122][4] , \row2_buffer[122][3] ,
         \row2_buffer[122][2] , \row2_buffer[122][1] , \row2_buffer[122][0] ,
         \row2_buffer[123][7] , \row2_buffer[123][6] , \row2_buffer[123][5] ,
         \row2_buffer[123][4] , \row2_buffer[123][3] , \row2_buffer[123][2] ,
         \row2_buffer[123][1] , \row2_buffer[123][0] , \row2_buffer[124][7] ,
         \row2_buffer[124][6] , \row2_buffer[124][5] , \row2_buffer[124][4] ,
         \row2_buffer[124][3] , \row2_buffer[124][2] , \row2_buffer[124][1] ,
         \row2_buffer[124][0] , \row2_buffer[125][7] , \row2_buffer[125][6] ,
         \row2_buffer[125][5] , \row2_buffer[125][4] , \row2_buffer[125][3] ,
         \row2_buffer[125][2] , \row2_buffer[125][1] , \row2_buffer[125][0] ,
         \row2_buffer[126][7] , \row2_buffer[126][6] , \row2_buffer[126][5] ,
         \row2_buffer[126][4] , \row2_buffer[126][3] , \row2_buffer[126][2] ,
         \row2_buffer[126][1] , \row2_buffer[126][0] , \row2_buffer[127][7] ,
         \row2_buffer[127][6] , \row2_buffer[127][5] , \row2_buffer[127][4] ,
         \row2_buffer[127][3] , \row2_buffer[127][2] , \row2_buffer[127][1] ,
         \row2_buffer[127][0] , \row2_buffer[128][7] , \row2_buffer[128][6] ,
         \row2_buffer[128][5] , \row2_buffer[128][4] , \row2_buffer[128][3] ,
         \row2_buffer[128][2] , \row2_buffer[128][1] , \row2_buffer[128][0] ,
         \row2_buffer[129][7] , \row2_buffer[129][6] , \row2_buffer[129][5] ,
         \row2_buffer[129][4] , \row2_buffer[129][3] , \row2_buffer[129][2] ,
         \row2_buffer[129][1] , \row2_buffer[129][0] , \row2_buffer[130][7] ,
         \row2_buffer[130][6] , \row2_buffer[130][5] , \row2_buffer[130][4] ,
         \row2_buffer[130][3] , \row2_buffer[130][2] , \row2_buffer[130][1] ,
         \row2_buffer[130][0] , \row2_buffer[131][7] , \row2_buffer[131][6] ,
         \row2_buffer[131][5] , \row2_buffer[131][4] , \row2_buffer[131][3] ,
         \row2_buffer[131][2] , \row2_buffer[131][1] , \row2_buffer[131][0] ,
         \row2_buffer[132][7] , \row2_buffer[132][6] , \row2_buffer[132][5] ,
         \row2_buffer[132][4] , \row2_buffer[132][3] , \row2_buffer[132][2] ,
         \row2_buffer[132][1] , \row2_buffer[132][0] , \row2_buffer[133][7] ,
         \row2_buffer[133][6] , \row2_buffer[133][5] , \row2_buffer[133][4] ,
         \row2_buffer[133][3] , \row2_buffer[133][2] , \row2_buffer[133][1] ,
         \row2_buffer[133][0] , \row2_buffer[134][7] , \row2_buffer[134][6] ,
         \row2_buffer[134][5] , \row2_buffer[134][4] , \row2_buffer[134][3] ,
         \row2_buffer[134][2] , \row2_buffer[134][1] , \row2_buffer[134][0] ,
         \row2_buffer[135][7] , \row2_buffer[135][6] , \row2_buffer[135][5] ,
         \row2_buffer[135][4] , \row2_buffer[135][3] , \row2_buffer[135][2] ,
         \row2_buffer[135][1] , \row2_buffer[135][0] , \row2_buffer[136][7] ,
         \row2_buffer[136][6] , \row2_buffer[136][5] , \row2_buffer[136][4] ,
         \row2_buffer[136][3] , \row2_buffer[136][2] , \row2_buffer[136][1] ,
         \row2_buffer[136][0] , \row2_buffer[137][7] , \row2_buffer[137][6] ,
         \row2_buffer[137][5] , \row2_buffer[137][4] , \row2_buffer[137][3] ,
         \row2_buffer[137][2] , \row2_buffer[137][1] , \row2_buffer[137][0] ,
         \row2_buffer[138][7] , \row2_buffer[138][6] , \row2_buffer[138][5] ,
         \row2_buffer[138][4] , \row2_buffer[138][3] , \row2_buffer[138][2] ,
         \row2_buffer[138][1] , \row2_buffer[138][0] , \row2_buffer[139][7] ,
         \row2_buffer[139][6] , \row2_buffer[139][5] , \row2_buffer[139][4] ,
         \row2_buffer[139][3] , \row2_buffer[139][2] , \row2_buffer[139][1] ,
         \row2_buffer[139][0] , \row2_buffer[140][7] , \row2_buffer[140][6] ,
         \row2_buffer[140][5] , \row2_buffer[140][4] , \row2_buffer[140][3] ,
         \row2_buffer[140][2] , \row2_buffer[140][1] , \row2_buffer[140][0] ,
         \row2_buffer[141][7] , \row2_buffer[141][6] , \row2_buffer[141][5] ,
         \row2_buffer[141][4] , \row2_buffer[141][3] , \row2_buffer[141][2] ,
         \row2_buffer[141][1] , \row2_buffer[141][0] , \row2_buffer[142][7] ,
         \row2_buffer[142][6] , \row2_buffer[142][5] , \row2_buffer[142][4] ,
         \row2_buffer[142][3] , \row2_buffer[142][2] , \row2_buffer[142][1] ,
         \row2_buffer[142][0] , \row2_buffer[143][7] , \row2_buffer[143][6] ,
         \row2_buffer[143][5] , \row2_buffer[143][4] , \row2_buffer[143][3] ,
         \row2_buffer[143][2] , \row2_buffer[143][1] , \row2_buffer[143][0] ,
         \row2_buffer[144][7] , \row2_buffer[144][6] , \row2_buffer[144][5] ,
         \row2_buffer[144][4] , \row2_buffer[144][3] , \row2_buffer[144][2] ,
         \row2_buffer[144][1] , \row2_buffer[144][0] , \row2_buffer[145][7] ,
         \row2_buffer[145][6] , \row2_buffer[145][5] , \row2_buffer[145][4] ,
         \row2_buffer[145][3] , \row2_buffer[145][2] , \row2_buffer[145][1] ,
         \row2_buffer[145][0] , \row2_buffer[146][7] , \row2_buffer[146][6] ,
         \row2_buffer[146][5] , \row2_buffer[146][4] , \row2_buffer[146][3] ,
         \row2_buffer[146][2] , \row2_buffer[146][1] , \row2_buffer[146][0] ,
         \row2_buffer[147][7] , \row2_buffer[147][6] , \row2_buffer[147][5] ,
         \row2_buffer[147][4] , \row2_buffer[147][3] , \row2_buffer[147][2] ,
         \row2_buffer[147][1] , \row2_buffer[147][0] , \row2_buffer[148][7] ,
         \row2_buffer[148][6] , \row2_buffer[148][5] , \row2_buffer[148][4] ,
         \row2_buffer[148][3] , \row2_buffer[148][2] , \row2_buffer[148][1] ,
         \row2_buffer[148][0] , \row2_buffer[149][7] , \row2_buffer[149][6] ,
         \row2_buffer[149][5] , \row2_buffer[149][4] , \row2_buffer[149][3] ,
         \row2_buffer[149][2] , \row2_buffer[149][1] , \row2_buffer[149][0] ,
         \row2_buffer[150][7] , \row2_buffer[150][6] , \row2_buffer[150][5] ,
         \row2_buffer[150][4] , \row2_buffer[150][3] , \row2_buffer[150][2] ,
         \row2_buffer[150][1] , \row2_buffer[150][0] , \row2_buffer[151][7] ,
         \row2_buffer[151][6] , \row2_buffer[151][5] , \row2_buffer[151][4] ,
         \row2_buffer[151][3] , \row2_buffer[151][2] , \row2_buffer[151][1] ,
         \row2_buffer[151][0] , \row2_buffer[152][7] , \row2_buffer[152][6] ,
         \row2_buffer[152][5] , \row2_buffer[152][4] , \row2_buffer[152][3] ,
         \row2_buffer[152][2] , \row2_buffer[152][1] , \row2_buffer[152][0] ,
         \row2_buffer[153][7] , \row2_buffer[153][6] , \row2_buffer[153][5] ,
         \row2_buffer[153][4] , \row2_buffer[153][3] , \row2_buffer[153][2] ,
         \row2_buffer[153][1] , \row2_buffer[153][0] , \row2_buffer[154][7] ,
         \row2_buffer[154][6] , \row2_buffer[154][5] , \row2_buffer[154][4] ,
         \row2_buffer[154][3] , \row2_buffer[154][2] , \row2_buffer[154][1] ,
         \row2_buffer[154][0] , \row2_buffer[155][7] , \row2_buffer[155][6] ,
         \row2_buffer[155][5] , \row2_buffer[155][4] , \row2_buffer[155][3] ,
         \row2_buffer[155][2] , \row2_buffer[155][1] , \row2_buffer[155][0] ,
         \row2_buffer[156][7] , \row2_buffer[156][6] , \row2_buffer[156][5] ,
         \row2_buffer[156][4] , \row2_buffer[156][3] , \row2_buffer[156][2] ,
         \row2_buffer[156][1] , \row2_buffer[156][0] , \row2_buffer[157][7] ,
         \row2_buffer[157][6] , \row2_buffer[157][5] , \row2_buffer[157][4] ,
         \row2_buffer[157][3] , \row2_buffer[157][2] , \row2_buffer[157][1] ,
         \row2_buffer[157][0] , \row2_buffer[158][7] , \row2_buffer[158][6] ,
         \row2_buffer[158][5] , \row2_buffer[158][4] , \row2_buffer[158][3] ,
         \row2_buffer[158][2] , \row2_buffer[158][1] , \row2_buffer[158][0] ,
         \row2_buffer[159][7] , \row2_buffer[159][6] , \row2_buffer[159][5] ,
         \row2_buffer[159][4] , \row2_buffer[159][3] , \row2_buffer[159][2] ,
         \row2_buffer[159][1] , \row2_buffer[159][0] , \row2_buffer[160][7] ,
         \row2_buffer[160][6] , \row2_buffer[160][5] , \row2_buffer[160][4] ,
         \row2_buffer[160][3] , \row2_buffer[160][2] , \row2_buffer[160][1] ,
         \row2_buffer[160][0] , \row2_buffer[161][7] , \row2_buffer[161][6] ,
         \row2_buffer[161][5] , \row2_buffer[161][4] , \row2_buffer[161][3] ,
         \row2_buffer[161][2] , \row2_buffer[161][1] , \row2_buffer[161][0] ,
         \row2_buffer[162][7] , \row2_buffer[162][6] , \row2_buffer[162][5] ,
         \row2_buffer[162][4] , \row2_buffer[162][3] , \row2_buffer[162][2] ,
         \row2_buffer[162][1] , \row2_buffer[162][0] , \row2_buffer[163][7] ,
         \row2_buffer[163][6] , \row2_buffer[163][5] , \row2_buffer[163][4] ,
         \row2_buffer[163][3] , \row2_buffer[163][2] , \row2_buffer[163][1] ,
         \row2_buffer[163][0] , \row2_buffer[164][7] , \row2_buffer[164][6] ,
         \row2_buffer[164][5] , \row2_buffer[164][4] , \row2_buffer[164][3] ,
         \row2_buffer[164][2] , \row2_buffer[164][1] , \row2_buffer[164][0] ,
         \row2_buffer[165][7] , \row2_buffer[165][6] , \row2_buffer[165][5] ,
         \row2_buffer[165][4] , \row2_buffer[165][3] , \row2_buffer[165][2] ,
         \row2_buffer[165][1] , \row2_buffer[165][0] , \row2_buffer[166][7] ,
         \row2_buffer[166][6] , \row2_buffer[166][5] , \row2_buffer[166][4] ,
         \row2_buffer[166][3] , \row2_buffer[166][2] , \row2_buffer[166][1] ,
         \row2_buffer[166][0] , \row2_buffer[167][7] , \row2_buffer[167][6] ,
         \row2_buffer[167][5] , \row2_buffer[167][4] , \row2_buffer[167][3] ,
         \row2_buffer[167][2] , \row2_buffer[167][1] , \row2_buffer[167][0] ,
         \row2_buffer[168][7] , \row2_buffer[168][6] , \row2_buffer[168][5] ,
         \row2_buffer[168][4] , \row2_buffer[168][3] , \row2_buffer[168][2] ,
         \row2_buffer[168][1] , \row2_buffer[168][0] , \row2_buffer[169][7] ,
         \row2_buffer[169][6] , \row2_buffer[169][5] , \row2_buffer[169][4] ,
         \row2_buffer[169][3] , \row2_buffer[169][2] , \row2_buffer[169][1] ,
         \row2_buffer[169][0] , \row2_buffer[170][7] , \row2_buffer[170][6] ,
         \row2_buffer[170][5] , \row2_buffer[170][4] , \row2_buffer[170][3] ,
         \row2_buffer[170][2] , \row2_buffer[170][1] , \row2_buffer[170][0] ,
         \row2_buffer[171][7] , \row2_buffer[171][6] , \row2_buffer[171][5] ,
         \row2_buffer[171][4] , \row2_buffer[171][3] , \row2_buffer[171][2] ,
         \row2_buffer[171][1] , \row2_buffer[171][0] , \row2_buffer[172][7] ,
         \row2_buffer[172][6] , \row2_buffer[172][5] , \row2_buffer[172][4] ,
         \row2_buffer[172][3] , \row2_buffer[172][2] , \row2_buffer[172][1] ,
         \row2_buffer[172][0] , \row2_buffer[173][7] , \row2_buffer[173][6] ,
         \row2_buffer[173][5] , \row2_buffer[173][4] , \row2_buffer[173][3] ,
         \row2_buffer[173][2] , \row2_buffer[173][1] , \row2_buffer[173][0] ,
         \row2_buffer[174][7] , \row2_buffer[174][6] , \row2_buffer[174][5] ,
         \row2_buffer[174][4] , \row2_buffer[174][3] , \row2_buffer[174][2] ,
         \row2_buffer[174][1] , \row2_buffer[174][0] , \row2_buffer[175][7] ,
         \row2_buffer[175][6] , \row2_buffer[175][5] , \row2_buffer[175][4] ,
         \row2_buffer[175][3] , \row2_buffer[175][2] , \row2_buffer[175][1] ,
         \row2_buffer[175][0] , \row2_buffer[176][7] , \row2_buffer[176][6] ,
         \row2_buffer[176][5] , \row2_buffer[176][4] , \row2_buffer[176][3] ,
         \row2_buffer[176][2] , \row2_buffer[176][1] , \row2_buffer[176][0] ,
         \row2_buffer[177][7] , \row2_buffer[177][6] , \row2_buffer[177][5] ,
         \row2_buffer[177][4] , \row2_buffer[177][3] , \row2_buffer[177][2] ,
         \row2_buffer[177][1] , \row2_buffer[177][0] , \row2_buffer[178][7] ,
         \row2_buffer[178][6] , \row2_buffer[178][5] , \row2_buffer[178][4] ,
         \row2_buffer[178][3] , \row2_buffer[178][2] , \row2_buffer[178][1] ,
         \row2_buffer[178][0] , \row2_buffer[179][7] , \row2_buffer[179][6] ,
         \row2_buffer[179][5] , \row2_buffer[179][4] , \row2_buffer[179][3] ,
         \row2_buffer[179][2] , \row2_buffer[179][1] , \row2_buffer[179][0] ,
         \row2_buffer[180][7] , \row2_buffer[180][6] , \row2_buffer[180][5] ,
         \row2_buffer[180][4] , \row2_buffer[180][3] , \row2_buffer[180][2] ,
         \row2_buffer[180][1] , \row2_buffer[180][0] , \row2_buffer[181][7] ,
         \row2_buffer[181][6] , \row2_buffer[181][5] , \row2_buffer[181][4] ,
         \row2_buffer[181][3] , \row2_buffer[181][2] , \row2_buffer[181][1] ,
         \row2_buffer[181][0] , \row2_buffer[182][7] , \row2_buffer[182][6] ,
         \row2_buffer[182][5] , \row2_buffer[182][4] , \row2_buffer[182][3] ,
         \row2_buffer[182][2] , \row2_buffer[182][1] , \row2_buffer[182][0] ,
         \row2_buffer[183][7] , \row2_buffer[183][6] , \row2_buffer[183][5] ,
         \row2_buffer[183][4] , \row2_buffer[183][3] , \row2_buffer[183][2] ,
         \row2_buffer[183][1] , \row2_buffer[183][0] , \row2_buffer[184][7] ,
         \row2_buffer[184][6] , \row2_buffer[184][5] , \row2_buffer[184][4] ,
         \row2_buffer[184][3] , \row2_buffer[184][2] , \row2_buffer[184][1] ,
         \row2_buffer[184][0] , \row2_buffer[185][7] , \row2_buffer[185][6] ,
         \row2_buffer[185][5] , \row2_buffer[185][4] , \row2_buffer[185][3] ,
         \row2_buffer[185][2] , \row2_buffer[185][1] , \row2_buffer[185][0] ,
         \row2_buffer[186][7] , \row2_buffer[186][6] , \row2_buffer[186][5] ,
         \row2_buffer[186][4] , \row2_buffer[186][3] , \row2_buffer[186][2] ,
         \row2_buffer[186][1] , \row2_buffer[186][0] , \row2_buffer[187][7] ,
         \row2_buffer[187][6] , \row2_buffer[187][5] , \row2_buffer[187][4] ,
         \row2_buffer[187][3] , \row2_buffer[187][2] , \row2_buffer[187][1] ,
         \row2_buffer[187][0] , \row2_buffer[188][7] , \row2_buffer[188][6] ,
         \row2_buffer[188][5] , \row2_buffer[188][4] , \row2_buffer[188][3] ,
         \row2_buffer[188][2] , \row2_buffer[188][1] , \row2_buffer[188][0] ,
         \row2_buffer[189][7] , \row2_buffer[189][6] , \row2_buffer[189][5] ,
         \row2_buffer[189][4] , \row2_buffer[189][3] , \row2_buffer[189][2] ,
         \row2_buffer[189][1] , \row2_buffer[189][0] , \row2_buffer[190][7] ,
         \row2_buffer[190][6] , \row2_buffer[190][5] , \row2_buffer[190][4] ,
         \row2_buffer[190][3] , \row2_buffer[190][2] , \row2_buffer[190][1] ,
         \row2_buffer[190][0] , \row2_buffer[191][7] , \row2_buffer[191][6] ,
         \row2_buffer[191][5] , \row2_buffer[191][4] , \row2_buffer[191][3] ,
         \row2_buffer[191][2] , \row2_buffer[191][1] , \row2_buffer[191][0] ,
         \row2_buffer[192][7] , \row2_buffer[192][6] , \row2_buffer[192][5] ,
         \row2_buffer[192][4] , \row2_buffer[192][3] , \row2_buffer[192][2] ,
         \row2_buffer[192][1] , \row2_buffer[192][0] , \row2_buffer[193][7] ,
         \row2_buffer[193][6] , \row2_buffer[193][5] , \row2_buffer[193][4] ,
         \row2_buffer[193][3] , \row2_buffer[193][2] , \row2_buffer[193][1] ,
         \row2_buffer[193][0] , \row2_buffer[194][7] , \row2_buffer[194][6] ,
         \row2_buffer[194][5] , \row2_buffer[194][4] , \row2_buffer[194][3] ,
         \row2_buffer[194][2] , \row2_buffer[194][1] , \row2_buffer[194][0] ,
         \row2_buffer[195][7] , \row2_buffer[195][6] , \row2_buffer[195][5] ,
         \row2_buffer[195][4] , \row2_buffer[195][3] , \row2_buffer[195][2] ,
         \row2_buffer[195][1] , \row2_buffer[195][0] , \row2_buffer[196][7] ,
         \row2_buffer[196][6] , \row2_buffer[196][5] , \row2_buffer[196][4] ,
         \row2_buffer[196][3] , \row2_buffer[196][2] , \row2_buffer[196][1] ,
         \row2_buffer[196][0] , \row2_buffer[197][7] , \row2_buffer[197][6] ,
         \row2_buffer[197][5] , \row2_buffer[197][4] , \row2_buffer[197][3] ,
         \row2_buffer[197][2] , \row2_buffer[197][1] , \row2_buffer[197][0] ,
         \row2_buffer[198][7] , \row2_buffer[198][6] , \row2_buffer[198][5] ,
         \row2_buffer[198][4] , \row2_buffer[198][3] , \row2_buffer[198][2] ,
         \row2_buffer[198][1] , \row2_buffer[198][0] , \row2_buffer[199][7] ,
         \row2_buffer[199][6] , \row2_buffer[199][5] , \row2_buffer[199][4] ,
         \row2_buffer[199][3] , \row2_buffer[199][2] , \row2_buffer[199][1] ,
         \row2_buffer[199][0] , \row2_buffer[200][7] , \row2_buffer[200][6] ,
         \row2_buffer[200][5] , \row2_buffer[200][4] , \row2_buffer[200][3] ,
         \row2_buffer[200][2] , \row2_buffer[200][1] , \row2_buffer[200][0] ,
         \row2_buffer[201][7] , \row2_buffer[201][6] , \row2_buffer[201][5] ,
         \row2_buffer[201][4] , \row2_buffer[201][3] , \row2_buffer[201][2] ,
         \row2_buffer[201][1] , \row2_buffer[201][0] , \row2_buffer[202][7] ,
         \row2_buffer[202][6] , \row2_buffer[202][5] , \row2_buffer[202][4] ,
         \row2_buffer[202][3] , \row2_buffer[202][2] , \row2_buffer[202][1] ,
         \row2_buffer[202][0] , \row2_buffer[203][7] , \row2_buffer[203][6] ,
         \row2_buffer[203][5] , \row2_buffer[203][4] , \row2_buffer[203][3] ,
         \row2_buffer[203][2] , \row2_buffer[203][1] , \row2_buffer[203][0] ,
         \row2_buffer[204][7] , \row2_buffer[204][6] , \row2_buffer[204][5] ,
         \row2_buffer[204][4] , \row2_buffer[204][3] , \row2_buffer[204][2] ,
         \row2_buffer[204][1] , \row2_buffer[204][0] , \row2_buffer[205][7] ,
         \row2_buffer[205][6] , \row2_buffer[205][5] , \row2_buffer[205][4] ,
         \row2_buffer[205][3] , \row2_buffer[205][2] , \row2_buffer[205][1] ,
         \row2_buffer[205][0] , \row2_buffer[206][7] , \row2_buffer[206][6] ,
         \row2_buffer[206][5] , \row2_buffer[206][4] , \row2_buffer[206][3] ,
         \row2_buffer[206][2] , \row2_buffer[206][1] , \row2_buffer[206][0] ,
         \row2_buffer[207][7] , \row2_buffer[207][6] , \row2_buffer[207][5] ,
         \row2_buffer[207][4] , \row2_buffer[207][3] , \row2_buffer[207][2] ,
         \row2_buffer[207][1] , \row2_buffer[207][0] , \row2_buffer[208][7] ,
         \row2_buffer[208][6] , \row2_buffer[208][5] , \row2_buffer[208][4] ,
         \row2_buffer[208][3] , \row2_buffer[208][2] , \row2_buffer[208][1] ,
         \row2_buffer[208][0] , \row2_buffer[209][7] , \row2_buffer[209][6] ,
         \row2_buffer[209][5] , \row2_buffer[209][4] , \row2_buffer[209][3] ,
         \row2_buffer[209][2] , \row2_buffer[209][1] , \row2_buffer[209][0] ,
         \row2_buffer[210][7] , \row2_buffer[210][6] , \row2_buffer[210][5] ,
         \row2_buffer[210][4] , \row2_buffer[210][3] , \row2_buffer[210][2] ,
         \row2_buffer[210][1] , \row2_buffer[210][0] , \row2_buffer[211][7] ,
         \row2_buffer[211][6] , \row2_buffer[211][5] , \row2_buffer[211][4] ,
         \row2_buffer[211][3] , \row2_buffer[211][2] , \row2_buffer[211][1] ,
         \row2_buffer[211][0] , \row2_buffer[212][7] , \row2_buffer[212][6] ,
         \row2_buffer[212][5] , \row2_buffer[212][4] , \row2_buffer[212][3] ,
         \row2_buffer[212][2] , \row2_buffer[212][1] , \row2_buffer[212][0] ,
         \row2_buffer[213][7] , \row2_buffer[213][6] , \row2_buffer[213][5] ,
         \row2_buffer[213][4] , \row2_buffer[213][3] , \row2_buffer[213][2] ,
         \row2_buffer[213][1] , \row2_buffer[213][0] , \row2_buffer[214][7] ,
         \row2_buffer[214][6] , \row2_buffer[214][5] , \row2_buffer[214][4] ,
         \row2_buffer[214][3] , \row2_buffer[214][2] , \row2_buffer[214][1] ,
         \row2_buffer[214][0] , \row2_buffer[215][7] , \row2_buffer[215][6] ,
         \row2_buffer[215][5] , \row2_buffer[215][4] , \row2_buffer[215][3] ,
         \row2_buffer[215][2] , \row2_buffer[215][1] , \row2_buffer[215][0] ,
         \row2_buffer[216][7] , \row2_buffer[216][6] , \row2_buffer[216][5] ,
         \row2_buffer[216][4] , \row2_buffer[216][3] , \row2_buffer[216][2] ,
         \row2_buffer[216][1] , \row2_buffer[216][0] , \row2_buffer[217][7] ,
         \row2_buffer[217][6] , \row2_buffer[217][5] , \row2_buffer[217][4] ,
         \row2_buffer[217][3] , \row2_buffer[217][2] , \row2_buffer[217][1] ,
         \row2_buffer[217][0] , \row2_buffer[218][7] , \row2_buffer[218][6] ,
         \row2_buffer[218][5] , \row2_buffer[218][4] , \row2_buffer[218][3] ,
         \row2_buffer[218][2] , \row2_buffer[218][1] , \row2_buffer[218][0] ,
         \row2_buffer[219][7] , \row2_buffer[219][6] , \row2_buffer[219][5] ,
         \row2_buffer[219][4] , \row2_buffer[219][3] , \row2_buffer[219][2] ,
         \row2_buffer[219][1] , \row2_buffer[219][0] , \row2_buffer[220][7] ,
         \row2_buffer[220][6] , \row2_buffer[220][5] , \row2_buffer[220][4] ,
         \row2_buffer[220][3] , \row2_buffer[220][2] , \row2_buffer[220][1] ,
         \row2_buffer[220][0] , \row2_buffer[221][7] , \row2_buffer[221][6] ,
         \row2_buffer[221][5] , \row2_buffer[221][4] , \row2_buffer[221][3] ,
         \row2_buffer[221][2] , \row2_buffer[221][1] , \row2_buffer[221][0] ,
         \row2_buffer[222][7] , \row2_buffer[222][6] , \row2_buffer[222][5] ,
         \row2_buffer[222][4] , \row2_buffer[222][3] , \row2_buffer[222][2] ,
         \row2_buffer[222][1] , \row2_buffer[222][0] , \row2_buffer[223][7] ,
         \row2_buffer[223][6] , \row2_buffer[223][5] , \row2_buffer[223][4] ,
         \row2_buffer[223][3] , \row2_buffer[223][2] , \row2_buffer[223][1] ,
         \row2_buffer[223][0] , \row2_buffer[224][7] , \row2_buffer[224][6] ,
         \row2_buffer[224][5] , \row2_buffer[224][4] , \row2_buffer[224][3] ,
         \row2_buffer[224][2] , \row2_buffer[224][1] , \row2_buffer[224][0] ,
         \row2_buffer[225][7] , \row2_buffer[225][6] , \row2_buffer[225][5] ,
         \row2_buffer[225][4] , \row2_buffer[225][3] , \row2_buffer[225][2] ,
         \row2_buffer[225][1] , \row2_buffer[225][0] , \row3_buffer[0][7] ,
         \row3_buffer[0][6] , \row3_buffer[0][5] , \row3_buffer[0][4] ,
         \row3_buffer[0][3] , \row3_buffer[0][2] , \row3_buffer[0][1] ,
         \row3_buffer[0][0] , \row3_buffer[1][7] , \row3_buffer[1][6] ,
         \row3_buffer[1][5] , \row3_buffer[1][4] , \row3_buffer[1][3] ,
         \row3_buffer[1][2] , \row3_buffer[1][1] , \row3_buffer[1][0] ,
         \row3_buffer[2][7] , \row3_buffer[2][6] , \row3_buffer[2][5] ,
         \row3_buffer[2][4] , \row3_buffer[2][3] , \row3_buffer[2][2] ,
         \row3_buffer[2][1] , \row3_buffer[2][0] , \row1_buffer[0][7] ,
         \row1_buffer[0][6] , \row1_buffer[0][5] , \row1_buffer[0][4] ,
         \row1_buffer[0][3] , \row1_buffer[0][2] , \row1_buffer[0][1] ,
         \row1_buffer[0][0] , \row1_buffer[1][7] , \row1_buffer[1][6] ,
         \row1_buffer[1][5] , \row1_buffer[1][4] , \row1_buffer[1][3] ,
         \row1_buffer[1][2] , \row1_buffer[1][1] , \row1_buffer[1][0] ,
         \row1_buffer[2][7] , \row1_buffer[2][6] , \row1_buffer[2][5] ,
         \row1_buffer[2][4] , \row1_buffer[2][3] , \row1_buffer[2][2] ,
         \row1_buffer[2][1] , \row1_buffer[2][0] , \row1_buffer[3][7] ,
         \row1_buffer[3][6] , \row1_buffer[3][5] , \row1_buffer[3][4] ,
         \row1_buffer[3][3] , \row1_buffer[3][2] , \row1_buffer[3][1] ,
         \row1_buffer[3][0] , \row1_buffer[4][7] , \row1_buffer[4][6] ,
         \row1_buffer[4][5] , \row1_buffer[4][4] , \row1_buffer[4][3] ,
         \row1_buffer[4][2] , \row1_buffer[4][1] , \row1_buffer[4][0] ,
         \row1_buffer[5][7] , \row1_buffer[5][6] , \row1_buffer[5][5] ,
         \row1_buffer[5][4] , \row1_buffer[5][3] , \row1_buffer[5][2] ,
         \row1_buffer[5][1] , \row1_buffer[5][0] , \row1_buffer[6][7] ,
         \row1_buffer[6][6] , \row1_buffer[6][5] , \row1_buffer[6][4] ,
         \row1_buffer[6][3] , \row1_buffer[6][2] , \row1_buffer[6][1] ,
         \row1_buffer[6][0] , \row1_buffer[7][7] , \row1_buffer[7][6] ,
         \row1_buffer[7][5] , \row1_buffer[7][4] , \row1_buffer[7][3] ,
         \row1_buffer[7][2] , \row1_buffer[7][1] , \row1_buffer[7][0] ,
         \row1_buffer[8][7] , \row1_buffer[8][6] , \row1_buffer[8][5] ,
         \row1_buffer[8][4] , \row1_buffer[8][3] , \row1_buffer[8][2] ,
         \row1_buffer[8][1] , \row1_buffer[8][0] , \row1_buffer[9][7] ,
         \row1_buffer[9][6] , \row1_buffer[9][5] , \row1_buffer[9][4] ,
         \row1_buffer[9][3] , \row1_buffer[9][2] , \row1_buffer[9][1] ,
         \row1_buffer[9][0] , \row1_buffer[10][7] , \row1_buffer[10][6] ,
         \row1_buffer[10][5] , \row1_buffer[10][4] , \row1_buffer[10][3] ,
         \row1_buffer[10][2] , \row1_buffer[10][1] , \row1_buffer[10][0] ,
         \row1_buffer[11][7] , \row1_buffer[11][6] , \row1_buffer[11][5] ,
         \row1_buffer[11][4] , \row1_buffer[11][3] , \row1_buffer[11][2] ,
         \row1_buffer[11][1] , \row1_buffer[11][0] , \row1_buffer[12][7] ,
         \row1_buffer[12][6] , \row1_buffer[12][5] , \row1_buffer[12][4] ,
         \row1_buffer[12][3] , \row1_buffer[12][2] , \row1_buffer[12][1] ,
         \row1_buffer[12][0] , \row1_buffer[13][7] , \row1_buffer[13][6] ,
         \row1_buffer[13][5] , \row1_buffer[13][4] , \row1_buffer[13][3] ,
         \row1_buffer[13][2] , \row1_buffer[13][1] , \row1_buffer[13][0] ,
         \row1_buffer[14][7] , \row1_buffer[14][6] , \row1_buffer[14][5] ,
         \row1_buffer[14][4] , \row1_buffer[14][3] , \row1_buffer[14][2] ,
         \row1_buffer[14][1] , \row1_buffer[14][0] , \row1_buffer[15][7] ,
         \row1_buffer[15][6] , \row1_buffer[15][5] , \row1_buffer[15][4] ,
         \row1_buffer[15][3] , \row1_buffer[15][2] , \row1_buffer[15][1] ,
         \row1_buffer[15][0] , \row1_buffer[16][7] , \row1_buffer[16][6] ,
         \row1_buffer[16][5] , \row1_buffer[16][4] , \row1_buffer[16][3] ,
         \row1_buffer[16][2] , \row1_buffer[16][1] , \row1_buffer[16][0] ,
         \row1_buffer[17][7] , \row1_buffer[17][6] , \row1_buffer[17][5] ,
         \row1_buffer[17][4] , \row1_buffer[17][3] , \row1_buffer[17][2] ,
         \row1_buffer[17][1] , \row1_buffer[17][0] , \row1_buffer[18][7] ,
         \row1_buffer[18][6] , \row1_buffer[18][5] , \row1_buffer[18][4] ,
         \row1_buffer[18][3] , \row1_buffer[18][2] , \row1_buffer[18][1] ,
         \row1_buffer[18][0] , \row1_buffer[19][7] , \row1_buffer[19][6] ,
         \row1_buffer[19][5] , \row1_buffer[19][4] , \row1_buffer[19][3] ,
         \row1_buffer[19][2] , \row1_buffer[19][1] , \row1_buffer[19][0] ,
         \row1_buffer[20][7] , \row1_buffer[20][6] , \row1_buffer[20][5] ,
         \row1_buffer[20][4] , \row1_buffer[20][3] , \row1_buffer[20][2] ,
         \row1_buffer[20][1] , \row1_buffer[20][0] , \row1_buffer[21][7] ,
         \row1_buffer[21][6] , \row1_buffer[21][5] , \row1_buffer[21][4] ,
         \row1_buffer[21][3] , \row1_buffer[21][2] , \row1_buffer[21][1] ,
         \row1_buffer[21][0] , \row1_buffer[22][7] , \row1_buffer[22][6] ,
         \row1_buffer[22][5] , \row1_buffer[22][4] , \row1_buffer[22][3] ,
         \row1_buffer[22][2] , \row1_buffer[22][1] , \row1_buffer[22][0] ,
         \row1_buffer[23][7] , \row1_buffer[23][6] , \row1_buffer[23][5] ,
         \row1_buffer[23][4] , \row1_buffer[23][3] , \row1_buffer[23][2] ,
         \row1_buffer[23][1] , \row1_buffer[23][0] , \row1_buffer[24][7] ,
         \row1_buffer[24][6] , \row1_buffer[24][5] , \row1_buffer[24][4] ,
         \row1_buffer[24][3] , \row1_buffer[24][2] , \row1_buffer[24][1] ,
         \row1_buffer[24][0] , \row1_buffer[25][7] , \row1_buffer[25][6] ,
         \row1_buffer[25][5] , \row1_buffer[25][4] , \row1_buffer[25][3] ,
         \row1_buffer[25][2] , \row1_buffer[25][1] , \row1_buffer[25][0] ,
         \row1_buffer[26][7] , \row1_buffer[26][6] , \row1_buffer[26][5] ,
         \row1_buffer[26][4] , \row1_buffer[26][3] , \row1_buffer[26][2] ,
         \row1_buffer[26][1] , \row1_buffer[26][0] , \row1_buffer[27][7] ,
         \row1_buffer[27][6] , \row1_buffer[27][5] , \row1_buffer[27][4] ,
         \row1_buffer[27][3] , \row1_buffer[27][2] , \row1_buffer[27][1] ,
         \row1_buffer[27][0] , \row1_buffer[28][7] , \row1_buffer[28][6] ,
         \row1_buffer[28][5] , \row1_buffer[28][4] , \row1_buffer[28][3] ,
         \row1_buffer[28][2] , \row1_buffer[28][1] , \row1_buffer[28][0] ,
         \row1_buffer[29][7] , \row1_buffer[29][6] , \row1_buffer[29][5] ,
         \row1_buffer[29][4] , \row1_buffer[29][3] , \row1_buffer[29][2] ,
         \row1_buffer[29][1] , \row1_buffer[29][0] , \row1_buffer[30][7] ,
         \row1_buffer[30][6] , \row1_buffer[30][5] , \row1_buffer[30][4] ,
         \row1_buffer[30][3] , \row1_buffer[30][2] , \row1_buffer[30][1] ,
         \row1_buffer[30][0] , \row1_buffer[31][7] , \row1_buffer[31][6] ,
         \row1_buffer[31][5] , \row1_buffer[31][4] , \row1_buffer[31][3] ,
         \row1_buffer[31][2] , \row1_buffer[31][1] , \row1_buffer[31][0] ,
         \row1_buffer[32][7] , \row1_buffer[32][6] , \row1_buffer[32][5] ,
         \row1_buffer[32][4] , \row1_buffer[32][3] , \row1_buffer[32][2] ,
         \row1_buffer[32][1] , \row1_buffer[32][0] , \row1_buffer[33][7] ,
         \row1_buffer[33][6] , \row1_buffer[33][5] , \row1_buffer[33][4] ,
         \row1_buffer[33][3] , \row1_buffer[33][2] , \row1_buffer[33][1] ,
         \row1_buffer[33][0] , \row1_buffer[34][7] , \row1_buffer[34][6] ,
         \row1_buffer[34][5] , \row1_buffer[34][4] , \row1_buffer[34][3] ,
         \row1_buffer[34][2] , \row1_buffer[34][1] , \row1_buffer[34][0] ,
         \row1_buffer[35][7] , \row1_buffer[35][6] , \row1_buffer[35][5] ,
         \row1_buffer[35][4] , \row1_buffer[35][3] , \row1_buffer[35][2] ,
         \row1_buffer[35][1] , \row1_buffer[35][0] , \row1_buffer[36][7] ,
         \row1_buffer[36][6] , \row1_buffer[36][5] , \row1_buffer[36][4] ,
         \row1_buffer[36][3] , \row1_buffer[36][2] , \row1_buffer[36][1] ,
         \row1_buffer[36][0] , \row1_buffer[37][7] , \row1_buffer[37][6] ,
         \row1_buffer[37][5] , \row1_buffer[37][4] , \row1_buffer[37][3] ,
         \row1_buffer[37][2] , \row1_buffer[37][1] , \row1_buffer[37][0] ,
         \row1_buffer[38][7] , \row1_buffer[38][6] , \row1_buffer[38][5] ,
         \row1_buffer[38][4] , \row1_buffer[38][3] , \row1_buffer[38][2] ,
         \row1_buffer[38][1] , \row1_buffer[38][0] , \row1_buffer[39][7] ,
         \row1_buffer[39][6] , \row1_buffer[39][5] , \row1_buffer[39][4] ,
         \row1_buffer[39][3] , \row1_buffer[39][2] , \row1_buffer[39][1] ,
         \row1_buffer[39][0] , \row1_buffer[40][7] , \row1_buffer[40][6] ,
         \row1_buffer[40][5] , \row1_buffer[40][4] , \row1_buffer[40][3] ,
         \row1_buffer[40][2] , \row1_buffer[40][1] , \row1_buffer[40][0] ,
         \row1_buffer[41][7] , \row1_buffer[41][6] , \row1_buffer[41][5] ,
         \row1_buffer[41][4] , \row1_buffer[41][3] , \row1_buffer[41][2] ,
         \row1_buffer[41][1] , \row1_buffer[41][0] , \row1_buffer[42][7] ,
         \row1_buffer[42][6] , \row1_buffer[42][5] , \row1_buffer[42][4] ,
         \row1_buffer[42][3] , \row1_buffer[42][2] , \row1_buffer[42][1] ,
         \row1_buffer[42][0] , \row1_buffer[43][7] , \row1_buffer[43][6] ,
         \row1_buffer[43][5] , \row1_buffer[43][4] , \row1_buffer[43][3] ,
         \row1_buffer[43][2] , \row1_buffer[43][1] , \row1_buffer[43][0] ,
         \row1_buffer[44][7] , \row1_buffer[44][6] , \row1_buffer[44][5] ,
         \row1_buffer[44][4] , \row1_buffer[44][3] , \row1_buffer[44][2] ,
         \row1_buffer[44][1] , \row1_buffer[44][0] , \row1_buffer[45][7] ,
         \row1_buffer[45][6] , \row1_buffer[45][5] , \row1_buffer[45][4] ,
         \row1_buffer[45][3] , \row1_buffer[45][2] , \row1_buffer[45][1] ,
         \row1_buffer[45][0] , \row1_buffer[46][7] , \row1_buffer[46][6] ,
         \row1_buffer[46][5] , \row1_buffer[46][4] , \row1_buffer[46][3] ,
         \row1_buffer[46][2] , \row1_buffer[46][1] , \row1_buffer[46][0] ,
         \row1_buffer[47][7] , \row1_buffer[47][6] , \row1_buffer[47][5] ,
         \row1_buffer[47][4] , \row1_buffer[47][3] , \row1_buffer[47][2] ,
         \row1_buffer[47][1] , \row1_buffer[47][0] , \row1_buffer[48][7] ,
         \row1_buffer[48][6] , \row1_buffer[48][5] , \row1_buffer[48][4] ,
         \row1_buffer[48][3] , \row1_buffer[48][2] , \row1_buffer[48][1] ,
         \row1_buffer[48][0] , \row1_buffer[49][7] , \row1_buffer[49][6] ,
         \row1_buffer[49][5] , \row1_buffer[49][4] , \row1_buffer[49][3] ,
         \row1_buffer[49][2] , \row1_buffer[49][1] , \row1_buffer[49][0] ,
         \row1_buffer[50][7] , \row1_buffer[50][6] , \row1_buffer[50][5] ,
         \row1_buffer[50][4] , \row1_buffer[50][3] , \row1_buffer[50][2] ,
         \row1_buffer[50][1] , \row1_buffer[50][0] , \row1_buffer[51][7] ,
         \row1_buffer[51][6] , \row1_buffer[51][5] , \row1_buffer[51][4] ,
         \row1_buffer[51][3] , \row1_buffer[51][2] , \row1_buffer[51][1] ,
         \row1_buffer[51][0] , \row1_buffer[52][7] , \row1_buffer[52][6] ,
         \row1_buffer[52][5] , \row1_buffer[52][4] , \row1_buffer[52][3] ,
         \row1_buffer[52][2] , \row1_buffer[52][1] , \row1_buffer[52][0] ,
         \row1_buffer[53][7] , \row1_buffer[53][6] , \row1_buffer[53][5] ,
         \row1_buffer[53][4] , \row1_buffer[53][3] , \row1_buffer[53][2] ,
         \row1_buffer[53][1] , \row1_buffer[53][0] , \row1_buffer[54][7] ,
         \row1_buffer[54][6] , \row1_buffer[54][5] , \row1_buffer[54][4] ,
         \row1_buffer[54][3] , \row1_buffer[54][2] , \row1_buffer[54][1] ,
         \row1_buffer[54][0] , \row1_buffer[55][7] , \row1_buffer[55][6] ,
         \row1_buffer[55][5] , \row1_buffer[55][4] , \row1_buffer[55][3] ,
         \row1_buffer[55][2] , \row1_buffer[55][1] , \row1_buffer[55][0] ,
         \row1_buffer[56][7] , \row1_buffer[56][6] , \row1_buffer[56][5] ,
         \row1_buffer[56][4] , \row1_buffer[56][3] , \row1_buffer[56][2] ,
         \row1_buffer[56][1] , \row1_buffer[56][0] , \row1_buffer[57][7] ,
         \row1_buffer[57][6] , \row1_buffer[57][5] , \row1_buffer[57][4] ,
         \row1_buffer[57][3] , \row1_buffer[57][2] , \row1_buffer[57][1] ,
         \row1_buffer[57][0] , \row1_buffer[58][7] , \row1_buffer[58][6] ,
         \row1_buffer[58][5] , \row1_buffer[58][4] , \row1_buffer[58][3] ,
         \row1_buffer[58][2] , \row1_buffer[58][1] , \row1_buffer[58][0] ,
         \row1_buffer[59][7] , \row1_buffer[59][6] , \row1_buffer[59][5] ,
         \row1_buffer[59][4] , \row1_buffer[59][3] , \row1_buffer[59][2] ,
         \row1_buffer[59][1] , \row1_buffer[59][0] , \row1_buffer[60][7] ,
         \row1_buffer[60][6] , \row1_buffer[60][5] , \row1_buffer[60][4] ,
         \row1_buffer[60][3] , \row1_buffer[60][2] , \row1_buffer[60][1] ,
         \row1_buffer[60][0] , \row1_buffer[61][7] , \row1_buffer[61][6] ,
         \row1_buffer[61][5] , \row1_buffer[61][4] , \row1_buffer[61][3] ,
         \row1_buffer[61][2] , \row1_buffer[61][1] , \row1_buffer[61][0] ,
         \row1_buffer[62][7] , \row1_buffer[62][6] , \row1_buffer[62][5] ,
         \row1_buffer[62][4] , \row1_buffer[62][3] , \row1_buffer[62][2] ,
         \row1_buffer[62][1] , \row1_buffer[62][0] , \row1_buffer[63][7] ,
         \row1_buffer[63][6] , \row1_buffer[63][5] , \row1_buffer[63][4] ,
         \row1_buffer[63][3] , \row1_buffer[63][2] , \row1_buffer[63][1] ,
         \row1_buffer[63][0] , \row1_buffer[64][7] , \row1_buffer[64][6] ,
         \row1_buffer[64][5] , \row1_buffer[64][4] , \row1_buffer[64][3] ,
         \row1_buffer[64][2] , \row1_buffer[64][1] , \row1_buffer[64][0] ,
         \row1_buffer[65][7] , \row1_buffer[65][6] , \row1_buffer[65][5] ,
         \row1_buffer[65][4] , \row1_buffer[65][3] , \row1_buffer[65][2] ,
         \row1_buffer[65][1] , \row1_buffer[65][0] , \row1_buffer[66][7] ,
         \row1_buffer[66][6] , \row1_buffer[66][5] , \row1_buffer[66][4] ,
         \row1_buffer[66][3] , \row1_buffer[66][2] , \row1_buffer[66][1] ,
         \row1_buffer[66][0] , \row1_buffer[67][7] , \row1_buffer[67][6] ,
         \row1_buffer[67][5] , \row1_buffer[67][4] , \row1_buffer[67][3] ,
         \row1_buffer[67][2] , \row1_buffer[67][1] , \row1_buffer[67][0] ,
         \row1_buffer[68][7] , \row1_buffer[68][6] , \row1_buffer[68][5] ,
         \row1_buffer[68][4] , \row1_buffer[68][3] , \row1_buffer[68][2] ,
         \row1_buffer[68][1] , \row1_buffer[68][0] , \row1_buffer[69][7] ,
         \row1_buffer[69][6] , \row1_buffer[69][5] , \row1_buffer[69][4] ,
         \row1_buffer[69][3] , \row1_buffer[69][2] , \row1_buffer[69][1] ,
         \row1_buffer[69][0] , \row1_buffer[70][7] , \row1_buffer[70][6] ,
         \row1_buffer[70][5] , \row1_buffer[70][4] , \row1_buffer[70][3] ,
         \row1_buffer[70][2] , \row1_buffer[70][1] , \row1_buffer[70][0] ,
         \row1_buffer[71][7] , \row1_buffer[71][6] , \row1_buffer[71][5] ,
         \row1_buffer[71][4] , \row1_buffer[71][3] , \row1_buffer[71][2] ,
         \row1_buffer[71][1] , \row1_buffer[71][0] , \row1_buffer[72][7] ,
         \row1_buffer[72][6] , \row1_buffer[72][5] , \row1_buffer[72][4] ,
         \row1_buffer[72][3] , \row1_buffer[72][2] , \row1_buffer[72][1] ,
         \row1_buffer[72][0] , \row1_buffer[73][7] , \row1_buffer[73][6] ,
         \row1_buffer[73][5] , \row1_buffer[73][4] , \row1_buffer[73][3] ,
         \row1_buffer[73][2] , \row1_buffer[73][1] , \row1_buffer[73][0] ,
         \row1_buffer[74][7] , \row1_buffer[74][6] , \row1_buffer[74][5] ,
         \row1_buffer[74][4] , \row1_buffer[74][3] , \row1_buffer[74][2] ,
         \row1_buffer[74][1] , \row1_buffer[74][0] , \row1_buffer[75][7] ,
         \row1_buffer[75][6] , \row1_buffer[75][5] , \row1_buffer[75][4] ,
         \row1_buffer[75][3] , \row1_buffer[75][2] , \row1_buffer[75][1] ,
         \row1_buffer[75][0] , \row1_buffer[76][7] , \row1_buffer[76][6] ,
         \row1_buffer[76][5] , \row1_buffer[76][4] , \row1_buffer[76][3] ,
         \row1_buffer[76][2] , \row1_buffer[76][1] , \row1_buffer[76][0] ,
         \row1_buffer[77][7] , \row1_buffer[77][6] , \row1_buffer[77][5] ,
         \row1_buffer[77][4] , \row1_buffer[77][3] , \row1_buffer[77][2] ,
         \row1_buffer[77][1] , \row1_buffer[77][0] , \row1_buffer[78][7] ,
         \row1_buffer[78][6] , \row1_buffer[78][5] , \row1_buffer[78][4] ,
         \row1_buffer[78][3] , \row1_buffer[78][2] , \row1_buffer[78][1] ,
         \row1_buffer[78][0] , \row1_buffer[79][7] , \row1_buffer[79][6] ,
         \row1_buffer[79][5] , \row1_buffer[79][4] , \row1_buffer[79][3] ,
         \row1_buffer[79][2] , \row1_buffer[79][1] , \row1_buffer[79][0] ,
         \row1_buffer[80][7] , \row1_buffer[80][6] , \row1_buffer[80][5] ,
         \row1_buffer[80][4] , \row1_buffer[80][3] , \row1_buffer[80][2] ,
         \row1_buffer[80][1] , \row1_buffer[80][0] , \row1_buffer[81][7] ,
         \row1_buffer[81][6] , \row1_buffer[81][5] , \row1_buffer[81][4] ,
         \row1_buffer[81][3] , \row1_buffer[81][2] , \row1_buffer[81][1] ,
         \row1_buffer[81][0] , \row1_buffer[82][7] , \row1_buffer[82][6] ,
         \row1_buffer[82][5] , \row1_buffer[82][4] , \row1_buffer[82][3] ,
         \row1_buffer[82][2] , \row1_buffer[82][1] , \row1_buffer[82][0] ,
         \row1_buffer[83][7] , \row1_buffer[83][6] , \row1_buffer[83][5] ,
         \row1_buffer[83][4] , \row1_buffer[83][3] , \row1_buffer[83][2] ,
         \row1_buffer[83][1] , \row1_buffer[83][0] , \row1_buffer[84][7] ,
         \row1_buffer[84][6] , \row1_buffer[84][5] , \row1_buffer[84][4] ,
         \row1_buffer[84][3] , \row1_buffer[84][2] , \row1_buffer[84][1] ,
         \row1_buffer[84][0] , \row1_buffer[85][7] , \row1_buffer[85][6] ,
         \row1_buffer[85][5] , \row1_buffer[85][4] , \row1_buffer[85][3] ,
         \row1_buffer[85][2] , \row1_buffer[85][1] , \row1_buffer[85][0] ,
         \row1_buffer[86][7] , \row1_buffer[86][6] , \row1_buffer[86][5] ,
         \row1_buffer[86][4] , \row1_buffer[86][3] , \row1_buffer[86][2] ,
         \row1_buffer[86][1] , \row1_buffer[86][0] , \row1_buffer[87][7] ,
         \row1_buffer[87][6] , \row1_buffer[87][5] , \row1_buffer[87][4] ,
         \row1_buffer[87][3] , \row1_buffer[87][2] , \row1_buffer[87][1] ,
         \row1_buffer[87][0] , \row1_buffer[88][7] , \row1_buffer[88][6] ,
         \row1_buffer[88][5] , \row1_buffer[88][4] , \row1_buffer[88][3] ,
         \row1_buffer[88][2] , \row1_buffer[88][1] , \row1_buffer[88][0] ,
         \row1_buffer[89][7] , \row1_buffer[89][6] , \row1_buffer[89][5] ,
         \row1_buffer[89][4] , \row1_buffer[89][3] , \row1_buffer[89][2] ,
         \row1_buffer[89][1] , \row1_buffer[89][0] , \row1_buffer[90][7] ,
         \row1_buffer[90][6] , \row1_buffer[90][5] , \row1_buffer[90][4] ,
         \row1_buffer[90][3] , \row1_buffer[90][2] , \row1_buffer[90][1] ,
         \row1_buffer[90][0] , \row1_buffer[91][7] , \row1_buffer[91][6] ,
         \row1_buffer[91][5] , \row1_buffer[91][4] , \row1_buffer[91][3] ,
         \row1_buffer[91][2] , \row1_buffer[91][1] , \row1_buffer[91][0] ,
         \row1_buffer[92][7] , \row1_buffer[92][6] , \row1_buffer[92][5] ,
         \row1_buffer[92][4] , \row1_buffer[92][3] , \row1_buffer[92][2] ,
         \row1_buffer[92][1] , \row1_buffer[92][0] , \row1_buffer[93][7] ,
         \row1_buffer[93][6] , \row1_buffer[93][5] , \row1_buffer[93][4] ,
         \row1_buffer[93][3] , \row1_buffer[93][2] , \row1_buffer[93][1] ,
         \row1_buffer[93][0] , \row1_buffer[94][7] , \row1_buffer[94][6] ,
         \row1_buffer[94][5] , \row1_buffer[94][4] , \row1_buffer[94][3] ,
         \row1_buffer[94][2] , \row1_buffer[94][1] , \row1_buffer[94][0] ,
         \row1_buffer[95][7] , \row1_buffer[95][6] , \row1_buffer[95][5] ,
         \row1_buffer[95][4] , \row1_buffer[95][3] , \row1_buffer[95][2] ,
         \row1_buffer[95][1] , \row1_buffer[95][0] , \row1_buffer[96][7] ,
         \row1_buffer[96][6] , \row1_buffer[96][5] , \row1_buffer[96][4] ,
         \row1_buffer[96][3] , \row1_buffer[96][2] , \row1_buffer[96][1] ,
         \row1_buffer[96][0] , \row1_buffer[97][7] , \row1_buffer[97][6] ,
         \row1_buffer[97][5] , \row1_buffer[97][4] , \row1_buffer[97][3] ,
         \row1_buffer[97][2] , \row1_buffer[97][1] , \row1_buffer[97][0] ,
         \row1_buffer[98][7] , \row1_buffer[98][6] , \row1_buffer[98][5] ,
         \row1_buffer[98][4] , \row1_buffer[98][3] , \row1_buffer[98][2] ,
         \row1_buffer[98][1] , \row1_buffer[98][0] , \row1_buffer[99][7] ,
         \row1_buffer[99][6] , \row1_buffer[99][5] , \row1_buffer[99][4] ,
         \row1_buffer[99][3] , \row1_buffer[99][2] , \row1_buffer[99][1] ,
         \row1_buffer[99][0] , \row1_buffer[100][7] , \row1_buffer[100][6] ,
         \row1_buffer[100][5] , \row1_buffer[100][4] , \row1_buffer[100][3] ,
         \row1_buffer[100][2] , \row1_buffer[100][1] , \row1_buffer[100][0] ,
         \row1_buffer[101][7] , \row1_buffer[101][6] , \row1_buffer[101][5] ,
         \row1_buffer[101][4] , \row1_buffer[101][3] , \row1_buffer[101][2] ,
         \row1_buffer[101][1] , \row1_buffer[101][0] , \row1_buffer[102][7] ,
         \row1_buffer[102][6] , \row1_buffer[102][5] , \row1_buffer[102][4] ,
         \row1_buffer[102][3] , \row1_buffer[102][2] , \row1_buffer[102][1] ,
         \row1_buffer[102][0] , \row1_buffer[103][7] , \row1_buffer[103][6] ,
         \row1_buffer[103][5] , \row1_buffer[103][4] , \row1_buffer[103][3] ,
         \row1_buffer[103][2] , \row1_buffer[103][1] , \row1_buffer[103][0] ,
         \row1_buffer[104][7] , \row1_buffer[104][6] , \row1_buffer[104][5] ,
         \row1_buffer[104][4] , \row1_buffer[104][3] , \row1_buffer[104][2] ,
         \row1_buffer[104][1] , \row1_buffer[104][0] , \row1_buffer[105][7] ,
         \row1_buffer[105][6] , \row1_buffer[105][5] , \row1_buffer[105][4] ,
         \row1_buffer[105][3] , \row1_buffer[105][2] , \row1_buffer[105][1] ,
         \row1_buffer[105][0] , \row1_buffer[106][7] , \row1_buffer[106][6] ,
         \row1_buffer[106][5] , \row1_buffer[106][4] , \row1_buffer[106][3] ,
         \row1_buffer[106][2] , \row1_buffer[106][1] , \row1_buffer[106][0] ,
         \row1_buffer[107][7] , \row1_buffer[107][6] , \row1_buffer[107][5] ,
         \row1_buffer[107][4] , \row1_buffer[107][3] , \row1_buffer[107][2] ,
         \row1_buffer[107][1] , \row1_buffer[107][0] , \row1_buffer[108][7] ,
         \row1_buffer[108][6] , \row1_buffer[108][5] , \row1_buffer[108][4] ,
         \row1_buffer[108][3] , \row1_buffer[108][2] , \row1_buffer[108][1] ,
         \row1_buffer[108][0] , \row1_buffer[109][7] , \row1_buffer[109][6] ,
         \row1_buffer[109][5] , \row1_buffer[109][4] , \row1_buffer[109][3] ,
         \row1_buffer[109][2] , \row1_buffer[109][1] , \row1_buffer[109][0] ,
         \row1_buffer[110][7] , \row1_buffer[110][6] , \row1_buffer[110][5] ,
         \row1_buffer[110][4] , \row1_buffer[110][3] , \row1_buffer[110][2] ,
         \row1_buffer[110][1] , \row1_buffer[110][0] , \row1_buffer[111][7] ,
         \row1_buffer[111][6] , \row1_buffer[111][5] , \row1_buffer[111][4] ,
         \row1_buffer[111][3] , \row1_buffer[111][2] , \row1_buffer[111][1] ,
         \row1_buffer[111][0] , \row1_buffer[112][7] , \row1_buffer[112][6] ,
         \row1_buffer[112][5] , \row1_buffer[112][4] , \row1_buffer[112][3] ,
         \row1_buffer[112][2] , \row1_buffer[112][1] , \row1_buffer[112][0] ,
         \row1_buffer[113][7] , \row1_buffer[113][6] , \row1_buffer[113][5] ,
         \row1_buffer[113][4] , \row1_buffer[113][3] , \row1_buffer[113][2] ,
         \row1_buffer[113][1] , \row1_buffer[113][0] , \row1_buffer[114][7] ,
         \row1_buffer[114][6] , \row1_buffer[114][5] , \row1_buffer[114][4] ,
         \row1_buffer[114][3] , \row1_buffer[114][2] , \row1_buffer[114][1] ,
         \row1_buffer[114][0] , \row1_buffer[115][7] , \row1_buffer[115][6] ,
         \row1_buffer[115][5] , \row1_buffer[115][4] , \row1_buffer[115][3] ,
         \row1_buffer[115][2] , \row1_buffer[115][1] , \row1_buffer[115][0] ,
         \row1_buffer[116][7] , \row1_buffer[116][6] , \row1_buffer[116][5] ,
         \row1_buffer[116][4] , \row1_buffer[116][3] , \row1_buffer[116][2] ,
         \row1_buffer[116][1] , \row1_buffer[116][0] , \row1_buffer[117][7] ,
         \row1_buffer[117][6] , \row1_buffer[117][5] , \row1_buffer[117][4] ,
         \row1_buffer[117][3] , \row1_buffer[117][2] , \row1_buffer[117][1] ,
         \row1_buffer[117][0] , \row1_buffer[118][7] , \row1_buffer[118][6] ,
         \row1_buffer[118][5] , \row1_buffer[118][4] , \row1_buffer[118][3] ,
         \row1_buffer[118][2] , \row1_buffer[118][1] , \row1_buffer[118][0] ,
         \row1_buffer[119][7] , \row1_buffer[119][6] , \row1_buffer[119][5] ,
         \row1_buffer[119][4] , \row1_buffer[119][3] , \row1_buffer[119][2] ,
         \row1_buffer[119][1] , \row1_buffer[119][0] , \row1_buffer[120][7] ,
         \row1_buffer[120][6] , \row1_buffer[120][5] , \row1_buffer[120][4] ,
         \row1_buffer[120][3] , \row1_buffer[120][2] , \row1_buffer[120][1] ,
         \row1_buffer[120][0] , \row1_buffer[121][7] , \row1_buffer[121][6] ,
         \row1_buffer[121][5] , \row1_buffer[121][4] , \row1_buffer[121][3] ,
         \row1_buffer[121][2] , \row1_buffer[121][1] , \row1_buffer[121][0] ,
         \row1_buffer[122][7] , \row1_buffer[122][6] , \row1_buffer[122][5] ,
         \row1_buffer[122][4] , \row1_buffer[122][3] , \row1_buffer[122][2] ,
         \row1_buffer[122][1] , \row1_buffer[122][0] , \row1_buffer[123][7] ,
         \row1_buffer[123][6] , \row1_buffer[123][5] , \row1_buffer[123][4] ,
         \row1_buffer[123][3] , \row1_buffer[123][2] , \row1_buffer[123][1] ,
         \row1_buffer[123][0] , \row1_buffer[124][7] , \row1_buffer[124][6] ,
         \row1_buffer[124][5] , \row1_buffer[124][4] , \row1_buffer[124][3] ,
         \row1_buffer[124][2] , \row1_buffer[124][1] , \row1_buffer[124][0] ,
         \row1_buffer[125][7] , \row1_buffer[125][6] , \row1_buffer[125][5] ,
         \row1_buffer[125][4] , \row1_buffer[125][3] , \row1_buffer[125][2] ,
         \row1_buffer[125][1] , \row1_buffer[125][0] , \row1_buffer[126][7] ,
         \row1_buffer[126][6] , \row1_buffer[126][5] , \row1_buffer[126][4] ,
         \row1_buffer[126][3] , \row1_buffer[126][2] , \row1_buffer[126][1] ,
         \row1_buffer[126][0] , \row1_buffer[127][7] , \row1_buffer[127][6] ,
         \row1_buffer[127][5] , \row1_buffer[127][4] , \row1_buffer[127][3] ,
         \row1_buffer[127][2] , \row1_buffer[127][1] , \row1_buffer[127][0] ,
         \row1_buffer[128][7] , \row1_buffer[128][6] , \row1_buffer[128][5] ,
         \row1_buffer[128][4] , \row1_buffer[128][3] , \row1_buffer[128][2] ,
         \row1_buffer[128][1] , \row1_buffer[128][0] , \row1_buffer[129][7] ,
         \row1_buffer[129][6] , \row1_buffer[129][5] , \row1_buffer[129][4] ,
         \row1_buffer[129][3] , \row1_buffer[129][2] , \row1_buffer[129][1] ,
         \row1_buffer[129][0] , \row1_buffer[130][7] , \row1_buffer[130][6] ,
         \row1_buffer[130][5] , \row1_buffer[130][4] , \row1_buffer[130][3] ,
         \row1_buffer[130][2] , \row1_buffer[130][1] , \row1_buffer[130][0] ,
         \row1_buffer[131][7] , \row1_buffer[131][6] , \row1_buffer[131][5] ,
         \row1_buffer[131][4] , \row1_buffer[131][3] , \row1_buffer[131][2] ,
         \row1_buffer[131][1] , \row1_buffer[131][0] , \row1_buffer[132][7] ,
         \row1_buffer[132][6] , \row1_buffer[132][5] , \row1_buffer[132][4] ,
         \row1_buffer[132][3] , \row1_buffer[132][2] , \row1_buffer[132][1] ,
         \row1_buffer[132][0] , \row1_buffer[133][7] , \row1_buffer[133][6] ,
         \row1_buffer[133][5] , \row1_buffer[133][4] , \row1_buffer[133][3] ,
         \row1_buffer[133][2] , \row1_buffer[133][1] , \row1_buffer[133][0] ,
         \row1_buffer[134][7] , \row1_buffer[134][6] , \row1_buffer[134][5] ,
         \row1_buffer[134][4] , \row1_buffer[134][3] , \row1_buffer[134][2] ,
         \row1_buffer[134][1] , \row1_buffer[134][0] , \row1_buffer[135][7] ,
         \row1_buffer[135][6] , \row1_buffer[135][5] , \row1_buffer[135][4] ,
         \row1_buffer[135][3] , \row1_buffer[135][2] , \row1_buffer[135][1] ,
         \row1_buffer[135][0] , \row1_buffer[136][7] , \row1_buffer[136][6] ,
         \row1_buffer[136][5] , \row1_buffer[136][4] , \row1_buffer[136][3] ,
         \row1_buffer[136][2] , \row1_buffer[136][1] , \row1_buffer[136][0] ,
         \row1_buffer[137][7] , \row1_buffer[137][6] , \row1_buffer[137][5] ,
         \row1_buffer[137][4] , \row1_buffer[137][3] , \row1_buffer[137][2] ,
         \row1_buffer[137][1] , \row1_buffer[137][0] , \row1_buffer[138][7] ,
         \row1_buffer[138][6] , \row1_buffer[138][5] , \row1_buffer[138][4] ,
         \row1_buffer[138][3] , \row1_buffer[138][2] , \row1_buffer[138][1] ,
         \row1_buffer[138][0] , \row1_buffer[139][7] , \row1_buffer[139][6] ,
         \row1_buffer[139][5] , \row1_buffer[139][4] , \row1_buffer[139][3] ,
         \row1_buffer[139][2] , \row1_buffer[139][1] , \row1_buffer[139][0] ,
         \row1_buffer[140][7] , \row1_buffer[140][6] , \row1_buffer[140][5] ,
         \row1_buffer[140][4] , \row1_buffer[140][3] , \row1_buffer[140][2] ,
         \row1_buffer[140][1] , \row1_buffer[140][0] , \row1_buffer[141][7] ,
         \row1_buffer[141][6] , \row1_buffer[141][5] , \row1_buffer[141][4] ,
         \row1_buffer[141][3] , \row1_buffer[141][2] , \row1_buffer[141][1] ,
         \row1_buffer[141][0] , \row1_buffer[142][7] , \row1_buffer[142][6] ,
         \row1_buffer[142][5] , \row1_buffer[142][4] , \row1_buffer[142][3] ,
         \row1_buffer[142][2] , \row1_buffer[142][1] , \row1_buffer[142][0] ,
         \row1_buffer[143][7] , \row1_buffer[143][6] , \row1_buffer[143][5] ,
         \row1_buffer[143][4] , \row1_buffer[143][3] , \row1_buffer[143][2] ,
         \row1_buffer[143][1] , \row1_buffer[143][0] , \row1_buffer[144][7] ,
         \row1_buffer[144][6] , \row1_buffer[144][5] , \row1_buffer[144][4] ,
         \row1_buffer[144][3] , \row1_buffer[144][2] , \row1_buffer[144][1] ,
         \row1_buffer[144][0] , \row1_buffer[145][7] , \row1_buffer[145][6] ,
         \row1_buffer[145][5] , \row1_buffer[145][4] , \row1_buffer[145][3] ,
         \row1_buffer[145][2] , \row1_buffer[145][1] , \row1_buffer[145][0] ,
         \row1_buffer[146][7] , \row1_buffer[146][6] , \row1_buffer[146][5] ,
         \row1_buffer[146][4] , \row1_buffer[146][3] , \row1_buffer[146][2] ,
         \row1_buffer[146][1] , \row1_buffer[146][0] , \row1_buffer[147][7] ,
         \row1_buffer[147][6] , \row1_buffer[147][5] , \row1_buffer[147][4] ,
         \row1_buffer[147][3] , \row1_buffer[147][2] , \row1_buffer[147][1] ,
         \row1_buffer[147][0] , \row1_buffer[148][7] , \row1_buffer[148][6] ,
         \row1_buffer[148][5] , \row1_buffer[148][4] , \row1_buffer[148][3] ,
         \row1_buffer[148][2] , \row1_buffer[148][1] , \row1_buffer[148][0] ,
         \row1_buffer[149][7] , \row1_buffer[149][6] , \row1_buffer[149][5] ,
         \row1_buffer[149][4] , \row1_buffer[149][3] , \row1_buffer[149][2] ,
         \row1_buffer[149][1] , \row1_buffer[149][0] , \row1_buffer[150][7] ,
         \row1_buffer[150][6] , \row1_buffer[150][5] , \row1_buffer[150][4] ,
         \row1_buffer[150][3] , \row1_buffer[150][2] , \row1_buffer[150][1] ,
         \row1_buffer[150][0] , \row1_buffer[151][7] , \row1_buffer[151][6] ,
         \row1_buffer[151][5] , \row1_buffer[151][4] , \row1_buffer[151][3] ,
         \row1_buffer[151][2] , \row1_buffer[151][1] , \row1_buffer[151][0] ,
         \row1_buffer[152][7] , \row1_buffer[152][6] , \row1_buffer[152][5] ,
         \row1_buffer[152][4] , \row1_buffer[152][3] , \row1_buffer[152][2] ,
         \row1_buffer[152][1] , \row1_buffer[152][0] , \row1_buffer[153][7] ,
         \row1_buffer[153][6] , \row1_buffer[153][5] , \row1_buffer[153][4] ,
         \row1_buffer[153][3] , \row1_buffer[153][2] , \row1_buffer[153][1] ,
         \row1_buffer[153][0] , \row1_buffer[154][7] , \row1_buffer[154][6] ,
         \row1_buffer[154][5] , \row1_buffer[154][4] , \row1_buffer[154][3] ,
         \row1_buffer[154][2] , \row1_buffer[154][1] , \row1_buffer[154][0] ,
         \row1_buffer[155][7] , \row1_buffer[155][6] , \row1_buffer[155][5] ,
         \row1_buffer[155][4] , \row1_buffer[155][3] , \row1_buffer[155][2] ,
         \row1_buffer[155][1] , \row1_buffer[155][0] , \row1_buffer[156][7] ,
         \row1_buffer[156][6] , \row1_buffer[156][5] , \row1_buffer[156][4] ,
         \row1_buffer[156][3] , \row1_buffer[156][2] , \row1_buffer[156][1] ,
         \row1_buffer[156][0] , \row1_buffer[157][7] , \row1_buffer[157][6] ,
         \row1_buffer[157][5] , \row1_buffer[157][4] , \row1_buffer[157][3] ,
         \row1_buffer[157][2] , \row1_buffer[157][1] , \row1_buffer[157][0] ,
         \row1_buffer[158][7] , \row1_buffer[158][6] , \row1_buffer[158][5] ,
         \row1_buffer[158][4] , \row1_buffer[158][3] , \row1_buffer[158][2] ,
         \row1_buffer[158][1] , \row1_buffer[158][0] , \row1_buffer[159][7] ,
         \row1_buffer[159][6] , \row1_buffer[159][5] , \row1_buffer[159][4] ,
         \row1_buffer[159][3] , \row1_buffer[159][2] , \row1_buffer[159][1] ,
         \row1_buffer[159][0] , \row1_buffer[160][7] , \row1_buffer[160][6] ,
         \row1_buffer[160][5] , \row1_buffer[160][4] , \row1_buffer[160][3] ,
         \row1_buffer[160][2] , \row1_buffer[160][1] , \row1_buffer[160][0] ,
         \row1_buffer[161][7] , \row1_buffer[161][6] , \row1_buffer[161][5] ,
         \row1_buffer[161][4] , \row1_buffer[161][3] , \row1_buffer[161][2] ,
         \row1_buffer[161][1] , \row1_buffer[161][0] , \row1_buffer[162][7] ,
         \row1_buffer[162][6] , \row1_buffer[162][5] , \row1_buffer[162][4] ,
         \row1_buffer[162][3] , \row1_buffer[162][2] , \row1_buffer[162][1] ,
         \row1_buffer[162][0] , \row1_buffer[163][7] , \row1_buffer[163][6] ,
         \row1_buffer[163][5] , \row1_buffer[163][4] , \row1_buffer[163][3] ,
         \row1_buffer[163][2] , \row1_buffer[163][1] , \row1_buffer[163][0] ,
         \row1_buffer[164][7] , \row1_buffer[164][6] , \row1_buffer[164][5] ,
         \row1_buffer[164][4] , \row1_buffer[164][3] , \row1_buffer[164][2] ,
         \row1_buffer[164][1] , \row1_buffer[164][0] , \row1_buffer[165][7] ,
         \row1_buffer[165][6] , \row1_buffer[165][5] , \row1_buffer[165][4] ,
         \row1_buffer[165][3] , \row1_buffer[165][2] , \row1_buffer[165][1] ,
         \row1_buffer[165][0] , \row1_buffer[166][7] , \row1_buffer[166][6] ,
         \row1_buffer[166][5] , \row1_buffer[166][4] , \row1_buffer[166][3] ,
         \row1_buffer[166][2] , \row1_buffer[166][1] , \row1_buffer[166][0] ,
         \row1_buffer[167][7] , \row1_buffer[167][6] , \row1_buffer[167][5] ,
         \row1_buffer[167][4] , \row1_buffer[167][3] , \row1_buffer[167][2] ,
         \row1_buffer[167][1] , \row1_buffer[167][0] , \row1_buffer[168][7] ,
         \row1_buffer[168][6] , \row1_buffer[168][5] , \row1_buffer[168][4] ,
         \row1_buffer[168][3] , \row1_buffer[168][2] , \row1_buffer[168][1] ,
         \row1_buffer[168][0] , \row1_buffer[169][7] , \row1_buffer[169][6] ,
         \row1_buffer[169][5] , \row1_buffer[169][4] , \row1_buffer[169][3] ,
         \row1_buffer[169][2] , \row1_buffer[169][1] , \row1_buffer[169][0] ,
         \row1_buffer[170][7] , \row1_buffer[170][6] , \row1_buffer[170][5] ,
         \row1_buffer[170][4] , \row1_buffer[170][3] , \row1_buffer[170][2] ,
         \row1_buffer[170][1] , \row1_buffer[170][0] , \row1_buffer[171][7] ,
         \row1_buffer[171][6] , \row1_buffer[171][5] , \row1_buffer[171][4] ,
         \row1_buffer[171][3] , \row1_buffer[171][2] , \row1_buffer[171][1] ,
         \row1_buffer[171][0] , \row1_buffer[172][7] , \row1_buffer[172][6] ,
         \row1_buffer[172][5] , \row1_buffer[172][4] , \row1_buffer[172][3] ,
         \row1_buffer[172][2] , \row1_buffer[172][1] , \row1_buffer[172][0] ,
         \row1_buffer[173][7] , \row1_buffer[173][6] , \row1_buffer[173][5] ,
         \row1_buffer[173][4] , \row1_buffer[173][3] , \row1_buffer[173][2] ,
         \row1_buffer[173][1] , \row1_buffer[173][0] , \row1_buffer[174][7] ,
         \row1_buffer[174][6] , \row1_buffer[174][5] , \row1_buffer[174][4] ,
         \row1_buffer[174][3] , \row1_buffer[174][2] , \row1_buffer[174][1] ,
         \row1_buffer[174][0] , \row1_buffer[175][7] , \row1_buffer[175][6] ,
         \row1_buffer[175][5] , \row1_buffer[175][4] , \row1_buffer[175][3] ,
         \row1_buffer[175][2] , \row1_buffer[175][1] , \row1_buffer[175][0] ,
         \row1_buffer[176][7] , \row1_buffer[176][6] , \row1_buffer[176][5] ,
         \row1_buffer[176][4] , \row1_buffer[176][3] , \row1_buffer[176][2] ,
         \row1_buffer[176][1] , \row1_buffer[176][0] , \row1_buffer[177][7] ,
         \row1_buffer[177][6] , \row1_buffer[177][5] , \row1_buffer[177][4] ,
         \row1_buffer[177][3] , \row1_buffer[177][2] , \row1_buffer[177][1] ,
         \row1_buffer[177][0] , \row1_buffer[178][7] , \row1_buffer[178][6] ,
         \row1_buffer[178][5] , \row1_buffer[178][4] , \row1_buffer[178][3] ,
         \row1_buffer[178][2] , \row1_buffer[178][1] , \row1_buffer[178][0] ,
         \row1_buffer[179][7] , \row1_buffer[179][6] , \row1_buffer[179][5] ,
         \row1_buffer[179][4] , \row1_buffer[179][3] , \row1_buffer[179][2] ,
         \row1_buffer[179][1] , \row1_buffer[179][0] , \row1_buffer[180][7] ,
         \row1_buffer[180][6] , \row1_buffer[180][5] , \row1_buffer[180][4] ,
         \row1_buffer[180][3] , \row1_buffer[180][2] , \row1_buffer[180][1] ,
         \row1_buffer[180][0] , \row1_buffer[181][7] , \row1_buffer[181][6] ,
         \row1_buffer[181][5] , \row1_buffer[181][4] , \row1_buffer[181][3] ,
         \row1_buffer[181][2] , \row1_buffer[181][1] , \row1_buffer[181][0] ,
         \row1_buffer[182][7] , \row1_buffer[182][6] , \row1_buffer[182][5] ,
         \row1_buffer[182][4] , \row1_buffer[182][3] , \row1_buffer[182][2] ,
         \row1_buffer[182][1] , \row1_buffer[182][0] , \row1_buffer[183][7] ,
         \row1_buffer[183][6] , \row1_buffer[183][5] , \row1_buffer[183][4] ,
         \row1_buffer[183][3] , \row1_buffer[183][2] , \row1_buffer[183][1] ,
         \row1_buffer[183][0] , \row1_buffer[184][7] , \row1_buffer[184][6] ,
         \row1_buffer[184][5] , \row1_buffer[184][4] , \row1_buffer[184][3] ,
         \row1_buffer[184][2] , \row1_buffer[184][1] , \row1_buffer[184][0] ,
         \row1_buffer[185][7] , \row1_buffer[185][6] , \row1_buffer[185][5] ,
         \row1_buffer[185][4] , \row1_buffer[185][3] , \row1_buffer[185][2] ,
         \row1_buffer[185][1] , \row1_buffer[185][0] , \row1_buffer[186][7] ,
         \row1_buffer[186][6] , \row1_buffer[186][5] , \row1_buffer[186][4] ,
         \row1_buffer[186][3] , \row1_buffer[186][2] , \row1_buffer[186][1] ,
         \row1_buffer[186][0] , \row1_buffer[187][7] , \row1_buffer[187][6] ,
         \row1_buffer[187][5] , \row1_buffer[187][4] , \row1_buffer[187][3] ,
         \row1_buffer[187][2] , \row1_buffer[187][1] , \row1_buffer[187][0] ,
         \row1_buffer[188][7] , \row1_buffer[188][6] , \row1_buffer[188][5] ,
         \row1_buffer[188][4] , \row1_buffer[188][3] , \row1_buffer[188][2] ,
         \row1_buffer[188][1] , \row1_buffer[188][0] , \row1_buffer[189][7] ,
         \row1_buffer[189][6] , \row1_buffer[189][5] , \row1_buffer[189][4] ,
         \row1_buffer[189][3] , \row1_buffer[189][2] , \row1_buffer[189][1] ,
         \row1_buffer[189][0] , \row1_buffer[190][7] , \row1_buffer[190][6] ,
         \row1_buffer[190][5] , \row1_buffer[190][4] , \row1_buffer[190][3] ,
         \row1_buffer[190][2] , \row1_buffer[190][1] , \row1_buffer[190][0] ,
         \row1_buffer[191][7] , \row1_buffer[191][6] , \row1_buffer[191][5] ,
         \row1_buffer[191][4] , \row1_buffer[191][3] , \row1_buffer[191][2] ,
         \row1_buffer[191][1] , \row1_buffer[191][0] , \row1_buffer[192][7] ,
         \row1_buffer[192][6] , \row1_buffer[192][5] , \row1_buffer[192][4] ,
         \row1_buffer[192][3] , \row1_buffer[192][2] , \row1_buffer[192][1] ,
         \row1_buffer[192][0] , \row1_buffer[193][7] , \row1_buffer[193][6] ,
         \row1_buffer[193][5] , \row1_buffer[193][4] , \row1_buffer[193][3] ,
         \row1_buffer[193][2] , \row1_buffer[193][1] , \row1_buffer[193][0] ,
         \row1_buffer[194][7] , \row1_buffer[194][6] , \row1_buffer[194][5] ,
         \row1_buffer[194][4] , \row1_buffer[194][3] , \row1_buffer[194][2] ,
         \row1_buffer[194][1] , \row1_buffer[194][0] , \row1_buffer[195][7] ,
         \row1_buffer[195][6] , \row1_buffer[195][5] , \row1_buffer[195][4] ,
         \row1_buffer[195][3] , \row1_buffer[195][2] , \row1_buffer[195][1] ,
         \row1_buffer[195][0] , \row1_buffer[196][7] , \row1_buffer[196][6] ,
         \row1_buffer[196][5] , \row1_buffer[196][4] , \row1_buffer[196][3] ,
         \row1_buffer[196][2] , \row1_buffer[196][1] , \row1_buffer[196][0] ,
         \row1_buffer[197][7] , \row1_buffer[197][6] , \row1_buffer[197][5] ,
         \row1_buffer[197][4] , \row1_buffer[197][3] , \row1_buffer[197][2] ,
         \row1_buffer[197][1] , \row1_buffer[197][0] , \row1_buffer[198][7] ,
         \row1_buffer[198][6] , \row1_buffer[198][5] , \row1_buffer[198][4] ,
         \row1_buffer[198][3] , \row1_buffer[198][2] , \row1_buffer[198][1] ,
         \row1_buffer[198][0] , \row1_buffer[199][7] , \row1_buffer[199][6] ,
         \row1_buffer[199][5] , \row1_buffer[199][4] , \row1_buffer[199][3] ,
         \row1_buffer[199][2] , \row1_buffer[199][1] , \row1_buffer[199][0] ,
         \row1_buffer[200][7] , \row1_buffer[200][6] , \row1_buffer[200][5] ,
         \row1_buffer[200][4] , \row1_buffer[200][3] , \row1_buffer[200][2] ,
         \row1_buffer[200][1] , \row1_buffer[200][0] , \row1_buffer[201][7] ,
         \row1_buffer[201][6] , \row1_buffer[201][5] , \row1_buffer[201][4] ,
         \row1_buffer[201][3] , \row1_buffer[201][2] , \row1_buffer[201][1] ,
         \row1_buffer[201][0] , \row1_buffer[202][7] , \row1_buffer[202][6] ,
         \row1_buffer[202][5] , \row1_buffer[202][4] , \row1_buffer[202][3] ,
         \row1_buffer[202][2] , \row1_buffer[202][1] , \row1_buffer[202][0] ,
         \row1_buffer[203][7] , \row1_buffer[203][6] , \row1_buffer[203][5] ,
         \row1_buffer[203][4] , \row1_buffer[203][3] , \row1_buffer[203][2] ,
         \row1_buffer[203][1] , \row1_buffer[203][0] , \row1_buffer[204][7] ,
         \row1_buffer[204][6] , \row1_buffer[204][5] , \row1_buffer[204][4] ,
         \row1_buffer[204][3] , \row1_buffer[204][2] , \row1_buffer[204][1] ,
         \row1_buffer[204][0] , \row1_buffer[205][7] , \row1_buffer[205][6] ,
         \row1_buffer[205][5] , \row1_buffer[205][4] , \row1_buffer[205][3] ,
         \row1_buffer[205][2] , \row1_buffer[205][1] , \row1_buffer[205][0] ,
         \row1_buffer[206][7] , \row1_buffer[206][6] , \row1_buffer[206][5] ,
         \row1_buffer[206][4] , \row1_buffer[206][3] , \row1_buffer[206][2] ,
         \row1_buffer[206][1] , \row1_buffer[206][0] , \row1_buffer[207][7] ,
         \row1_buffer[207][6] , \row1_buffer[207][5] , \row1_buffer[207][4] ,
         \row1_buffer[207][3] , \row1_buffer[207][2] , \row1_buffer[207][1] ,
         \row1_buffer[207][0] , \row1_buffer[208][7] , \row1_buffer[208][6] ,
         \row1_buffer[208][5] , \row1_buffer[208][4] , \row1_buffer[208][3] ,
         \row1_buffer[208][2] , \row1_buffer[208][1] , \row1_buffer[208][0] ,
         \row1_buffer[209][7] , \row1_buffer[209][6] , \row1_buffer[209][5] ,
         \row1_buffer[209][4] , \row1_buffer[209][3] , \row1_buffer[209][2] ,
         \row1_buffer[209][1] , \row1_buffer[209][0] , \row1_buffer[210][7] ,
         \row1_buffer[210][6] , \row1_buffer[210][5] , \row1_buffer[210][4] ,
         \row1_buffer[210][3] , \row1_buffer[210][2] , \row1_buffer[210][1] ,
         \row1_buffer[210][0] , \row1_buffer[211][7] , \row1_buffer[211][6] ,
         \row1_buffer[211][5] , \row1_buffer[211][4] , \row1_buffer[211][3] ,
         \row1_buffer[211][2] , \row1_buffer[211][1] , \row1_buffer[211][0] ,
         \row1_buffer[212][7] , \row1_buffer[212][6] , \row1_buffer[212][5] ,
         \row1_buffer[212][4] , \row1_buffer[212][3] , \row1_buffer[212][2] ,
         \row1_buffer[212][1] , \row1_buffer[212][0] , \row1_buffer[213][7] ,
         \row1_buffer[213][6] , \row1_buffer[213][5] , \row1_buffer[213][4] ,
         \row1_buffer[213][3] , \row1_buffer[213][2] , \row1_buffer[213][1] ,
         \row1_buffer[213][0] , \row1_buffer[214][7] , \row1_buffer[214][6] ,
         \row1_buffer[214][5] , \row1_buffer[214][4] , \row1_buffer[214][3] ,
         \row1_buffer[214][2] , \row1_buffer[214][1] , \row1_buffer[214][0] ,
         \row1_buffer[215][7] , \row1_buffer[215][6] , \row1_buffer[215][5] ,
         \row1_buffer[215][4] , \row1_buffer[215][3] , \row1_buffer[215][2] ,
         \row1_buffer[215][1] , \row1_buffer[215][0] , \row1_buffer[216][7] ,
         \row1_buffer[216][6] , \row1_buffer[216][5] , \row1_buffer[216][4] ,
         \row1_buffer[216][3] , \row1_buffer[216][2] , \row1_buffer[216][1] ,
         \row1_buffer[216][0] , \row1_buffer[217][7] , \row1_buffer[217][6] ,
         \row1_buffer[217][5] , \row1_buffer[217][4] , \row1_buffer[217][3] ,
         \row1_buffer[217][2] , \row1_buffer[217][1] , \row1_buffer[217][0] ,
         \row1_buffer[218][7] , \row1_buffer[218][6] , \row1_buffer[218][5] ,
         \row1_buffer[218][4] , \row1_buffer[218][3] , \row1_buffer[218][2] ,
         \row1_buffer[218][1] , \row1_buffer[218][0] , \row1_buffer[219][7] ,
         \row1_buffer[219][6] , \row1_buffer[219][5] , \row1_buffer[219][4] ,
         \row1_buffer[219][3] , \row1_buffer[219][2] , \row1_buffer[219][1] ,
         \row1_buffer[219][0] , \row1_buffer[220][7] , \row1_buffer[220][6] ,
         \row1_buffer[220][5] , \row1_buffer[220][4] , \row1_buffer[220][3] ,
         \row1_buffer[220][2] , \row1_buffer[220][1] , \row1_buffer[220][0] ,
         \row1_buffer[221][7] , \row1_buffer[221][6] , \row1_buffer[221][5] ,
         \row1_buffer[221][4] , \row1_buffer[221][3] , \row1_buffer[221][2] ,
         \row1_buffer[221][1] , \row1_buffer[221][0] , \row1_buffer[222][7] ,
         \row1_buffer[222][6] , \row1_buffer[222][5] , \row1_buffer[222][4] ,
         \row1_buffer[222][3] , \row1_buffer[222][2] , \row1_buffer[222][1] ,
         \row1_buffer[222][0] , \row1_buffer[223][7] , \row1_buffer[223][6] ,
         \row1_buffer[223][5] , \row1_buffer[223][4] , \row1_buffer[223][3] ,
         \row1_buffer[223][2] , \row1_buffer[223][1] , \row1_buffer[223][0] ,
         \row1_buffer[224][7] , \row1_buffer[224][6] , \row1_buffer[224][5] ,
         \row1_buffer[224][4] , \row1_buffer[224][3] , \row1_buffer[224][2] ,
         \row1_buffer[224][1] , \row1_buffer[224][0] , \row1_buffer[225][7] ,
         \row1_buffer[225][6] , \row1_buffer[225][5] , \row1_buffer[225][4] ,
         \row1_buffer[225][3] , \row1_buffer[225][2] , \row1_buffer[225][1] ,
         \row1_buffer[225][0] ;

  DFFQX2 \pixel_22_reg[6]  ( .D(\row3_buffer[2][6] ), .CK(clk), .Q(pixel_22[6]) );
  DFFQX2 \pixel_21_reg[6]  ( .D(\row3_buffer[1][6] ), .CK(clk), .Q(pixel_21[6]) );
  DFFQX2 \pixel_20_reg[6]  ( .D(\row3_buffer[0][6] ), .CK(clk), .Q(pixel_20[6]) );
  DFFQX2 \pixel_12_reg[6]  ( .D(\row2_buffer[2][6] ), .CK(clk), .Q(pixel_12[6]) );
  DFFQX2 \pixel_11_reg[6]  ( .D(\row2_buffer[1][6] ), .CK(clk), .Q(pixel_11[6]) );
  DFFQX2 \pixel_10_reg[6]  ( .D(\row2_buffer[0][6] ), .CK(clk), .Q(pixel_10[6]) );
  DFFQX2 \pixel_02_reg[6]  ( .D(\row1_buffer[2][6] ), .CK(clk), .Q(pixel_02[6]) );
  DFFQX2 \pixel_00_reg[6]  ( .D(\row1_buffer[0][6] ), .CK(clk), .Q(pixel_00[6]) );
  DFFQX2 \pixel_01_reg[6]  ( .D(\row1_buffer[1][6] ), .CK(clk), .Q(pixel_01[6]) );
  DFFQXL \pixel_22_reg[7]  ( .D(\row3_buffer[2][7] ), .CK(clk), .Q(pixel_22[7]) );
  DFFQXL \pixel_21_reg[7]  ( .D(\row3_buffer[1][7] ), .CK(clk), .Q(pixel_21[7]) );
  DFFQXL \pixel_20_reg[7]  ( .D(\row3_buffer[0][7] ), .CK(clk), .Q(pixel_20[7]) );
  DFFQXL \pixel_12_reg[7]  ( .D(\row2_buffer[2][7] ), .CK(clk), .Q(pixel_12[7]) );
  DFFQXL \pixel_11_reg[7]  ( .D(\row2_buffer[1][7] ), .CK(clk), .Q(pixel_11[7]) );
  DFFQXL \pixel_10_reg[7]  ( .D(\row2_buffer[0][7] ), .CK(clk), .Q(pixel_10[7]) );
  DFFQXL \pixel_02_reg[7]  ( .D(\row1_buffer[2][7] ), .CK(clk), .Q(pixel_02[7]) );
  DFFQXL \pixel_00_reg[7]  ( .D(\row1_buffer[0][7] ), .CK(clk), .Q(pixel_00[7]) );
  DFFQXL \pixel_01_reg[7]  ( .D(\row1_buffer[1][7] ), .CK(clk), .Q(pixel_01[7]) );
  DFFQX2 \pixel_22_reg[0]  ( .D(\row3_buffer[2][0] ), .CK(clk), .Q(pixel_22[0]) );
  DFFQX2 \pixel_21_reg[0]  ( .D(\row3_buffer[1][0] ), .CK(clk), .Q(pixel_21[0]) );
  DFFQX2 \pixel_20_reg[0]  ( .D(\row3_buffer[0][0] ), .CK(clk), .Q(pixel_20[0]) );
  DFFQX2 \pixel_12_reg[0]  ( .D(\row2_buffer[2][0] ), .CK(clk), .Q(pixel_12[0]) );
  DFFQX2 \pixel_11_reg[0]  ( .D(\row2_buffer[1][0] ), .CK(clk), .Q(pixel_11[0]) );
  DFFQX2 \pixel_10_reg[0]  ( .D(\row2_buffer[0][0] ), .CK(clk), .Q(pixel_10[0]) );
  DFFQX2 \pixel_02_reg[0]  ( .D(\row1_buffer[2][0] ), .CK(clk), .Q(pixel_02[0]) );
  DFFQX2 \pixel_00_reg[0]  ( .D(\row1_buffer[0][0] ), .CK(clk), .Q(pixel_00[0]) );
  DFFQX2 \pixel_01_reg[0]  ( .D(\row1_buffer[1][0] ), .CK(clk), .Q(pixel_01[0]) );
  DFFQX2 \pixel_22_reg[4]  ( .D(\row3_buffer[2][4] ), .CK(clk), .Q(pixel_22[4]) );
  DFFQX2 \pixel_21_reg[4]  ( .D(\row3_buffer[1][4] ), .CK(clk), .Q(pixel_21[4]) );
  DFFQX2 \pixel_20_reg[4]  ( .D(\row3_buffer[0][4] ), .CK(clk), .Q(pixel_20[4]) );
  DFFQX2 \pixel_12_reg[4]  ( .D(\row2_buffer[2][4] ), .CK(clk), .Q(pixel_12[4]) );
  DFFQX2 \pixel_11_reg[4]  ( .D(\row2_buffer[1][4] ), .CK(clk), .Q(pixel_11[4]) );
  DFFQX2 \pixel_10_reg[4]  ( .D(\row2_buffer[0][4] ), .CK(clk), .Q(pixel_10[4]) );
  DFFQX2 \pixel_02_reg[4]  ( .D(\row1_buffer[2][4] ), .CK(clk), .Q(pixel_02[4]) );
  DFFQX2 \pixel_22_reg[2]  ( .D(\row3_buffer[2][2] ), .CK(clk), .Q(pixel_22[2]) );
  DFFQX2 \pixel_21_reg[2]  ( .D(\row3_buffer[1][2] ), .CK(clk), .Q(pixel_21[2]) );
  DFFQX2 \pixel_20_reg[2]  ( .D(\row3_buffer[0][2] ), .CK(clk), .Q(pixel_20[2]) );
  DFFQX2 \pixel_12_reg[2]  ( .D(\row2_buffer[2][2] ), .CK(clk), .Q(pixel_12[2]) );
  DFFQX2 \pixel_11_reg[2]  ( .D(\row2_buffer[1][2] ), .CK(clk), .Q(pixel_11[2]) );
  DFFQX2 \pixel_10_reg[2]  ( .D(\row2_buffer[0][2] ), .CK(clk), .Q(pixel_10[2]) );
  DFFQX2 \pixel_02_reg[2]  ( .D(\row1_buffer[2][2] ), .CK(clk), .Q(pixel_02[2]) );
  DFFQX2 \pixel_00_reg[4]  ( .D(\row1_buffer[0][4] ), .CK(clk), .Q(pixel_00[4]) );
  DFFQX2 \pixel_00_reg[2]  ( .D(\row1_buffer[0][2] ), .CK(clk), .Q(pixel_00[2]) );
  DFFQX2 \pixel_01_reg[4]  ( .D(\row1_buffer[1][4] ), .CK(clk), .Q(pixel_01[4]) );
  DFFQX2 \pixel_01_reg[2]  ( .D(\row1_buffer[1][2] ), .CK(clk), .Q(pixel_01[2]) );
  DFFQX2 \pixel_22_reg[1]  ( .D(\row3_buffer[2][1] ), .CK(clk), .Q(pixel_22[1]) );
  DFFQX2 \pixel_21_reg[1]  ( .D(\row3_buffer[1][1] ), .CK(clk), .Q(pixel_21[1]) );
  DFFQX2 \pixel_20_reg[1]  ( .D(\row3_buffer[0][1] ), .CK(clk), .Q(pixel_20[1]) );
  DFFQX2 \pixel_12_reg[1]  ( .D(\row2_buffer[2][1] ), .CK(clk), .Q(pixel_12[1]) );
  DFFQX2 \pixel_11_reg[1]  ( .D(\row2_buffer[1][1] ), .CK(clk), .Q(pixel_11[1]) );
  DFFQX2 \pixel_10_reg[1]  ( .D(\row2_buffer[0][1] ), .CK(clk), .Q(pixel_10[1]) );
  DFFQX2 \pixel_02_reg[1]  ( .D(\row1_buffer[2][1] ), .CK(clk), .Q(pixel_02[1]) );
  DFFQX2 \pixel_00_reg[1]  ( .D(\row1_buffer[0][1] ), .CK(clk), .Q(pixel_00[1]) );
  DFFQX2 \pixel_01_reg[1]  ( .D(\row1_buffer[1][1] ), .CK(clk), .Q(pixel_01[1]) );
  DFFQXL \row1_buffer_reg[0][6]  ( .D(\row1_buffer[1][6] ), .CK(clk), .Q(
        \row1_buffer[0][6] ) );
  DFFQXL \row1_buffer_reg[0][4]  ( .D(\row1_buffer[1][4] ), .CK(clk), .Q(
        \row1_buffer[0][4] ) );
  DFFQXL \row1_buffer_reg[0][2]  ( .D(\row1_buffer[1][2] ), .CK(clk), .Q(
        \row1_buffer[0][2] ) );
  DFFQXL \row1_buffer_reg[0][1]  ( .D(\row1_buffer[1][1] ), .CK(clk), .Q(
        \row1_buffer[0][1] ) );
  DFFQXL \row1_buffer_reg[0][0]  ( .D(\row1_buffer[1][0] ), .CK(clk), .Q(
        \row1_buffer[0][0] ) );
  DFFQXL \row1_buffer_reg[0][7]  ( .D(\row1_buffer[1][7] ), .CK(clk), .Q(
        \row1_buffer[0][7] ) );
  DFFQXL \row2_buffer_reg[225][7]  ( .D(\row3_buffer[0][7] ), .CK(clk), .Q(
        \row2_buffer[225][7] ) );
  DFFQXL \row2_buffer_reg[224][7]  ( .D(\row2_buffer[225][7] ), .CK(clk), .Q(
        \row2_buffer[224][7] ) );
  DFFQXL \row2_buffer_reg[223][7]  ( .D(\row2_buffer[224][7] ), .CK(clk), .Q(
        \row2_buffer[223][7] ) );
  DFFQXL \row2_buffer_reg[222][7]  ( .D(\row2_buffer[223][7] ), .CK(clk), .Q(
        \row2_buffer[222][7] ) );
  DFFQXL \row2_buffer_reg[221][7]  ( .D(\row2_buffer[222][7] ), .CK(clk), .Q(
        \row2_buffer[221][7] ) );
  DFFQXL \row2_buffer_reg[220][7]  ( .D(\row2_buffer[221][7] ), .CK(clk), .Q(
        \row2_buffer[220][7] ) );
  DFFQXL \row2_buffer_reg[219][7]  ( .D(\row2_buffer[220][7] ), .CK(clk), .Q(
        \row2_buffer[219][7] ) );
  DFFQXL \row2_buffer_reg[218][7]  ( .D(\row2_buffer[219][7] ), .CK(clk), .Q(
        \row2_buffer[218][7] ) );
  DFFQXL \row2_buffer_reg[217][7]  ( .D(\row2_buffer[218][7] ), .CK(clk), .Q(
        \row2_buffer[217][7] ) );
  DFFQXL \row2_buffer_reg[216][7]  ( .D(\row2_buffer[217][7] ), .CK(clk), .Q(
        \row2_buffer[216][7] ) );
  DFFQXL \row2_buffer_reg[215][7]  ( .D(\row2_buffer[216][7] ), .CK(clk), .Q(
        \row2_buffer[215][7] ) );
  DFFQXL \row2_buffer_reg[214][7]  ( .D(\row2_buffer[215][7] ), .CK(clk), .Q(
        \row2_buffer[214][7] ) );
  DFFQXL \row2_buffer_reg[213][7]  ( .D(\row2_buffer[214][7] ), .CK(clk), .Q(
        \row2_buffer[213][7] ) );
  DFFQXL \row2_buffer_reg[212][7]  ( .D(\row2_buffer[213][7] ), .CK(clk), .Q(
        \row2_buffer[212][7] ) );
  DFFQXL \row2_buffer_reg[211][7]  ( .D(\row2_buffer[212][7] ), .CK(clk), .Q(
        \row2_buffer[211][7] ) );
  DFFQXL \row2_buffer_reg[210][7]  ( .D(\row2_buffer[211][7] ), .CK(clk), .Q(
        \row2_buffer[210][7] ) );
  DFFQXL \row2_buffer_reg[209][7]  ( .D(\row2_buffer[210][7] ), .CK(clk), .Q(
        \row2_buffer[209][7] ) );
  DFFQXL \row2_buffer_reg[208][7]  ( .D(\row2_buffer[209][7] ), .CK(clk), .Q(
        \row2_buffer[208][7] ) );
  DFFQXL \row2_buffer_reg[207][7]  ( .D(\row2_buffer[208][7] ), .CK(clk), .Q(
        \row2_buffer[207][7] ) );
  DFFQXL \row2_buffer_reg[206][7]  ( .D(\row2_buffer[207][7] ), .CK(clk), .Q(
        \row2_buffer[206][7] ) );
  DFFQXL \row2_buffer_reg[205][7]  ( .D(\row2_buffer[206][7] ), .CK(clk), .Q(
        \row2_buffer[205][7] ) );
  DFFQXL \row2_buffer_reg[204][7]  ( .D(\row2_buffer[205][7] ), .CK(clk), .Q(
        \row2_buffer[204][7] ) );
  DFFQXL \row2_buffer_reg[203][7]  ( .D(\row2_buffer[204][7] ), .CK(clk), .Q(
        \row2_buffer[203][7] ) );
  DFFQXL \row2_buffer_reg[202][7]  ( .D(\row2_buffer[203][7] ), .CK(clk), .Q(
        \row2_buffer[202][7] ) );
  DFFQXL \row2_buffer_reg[201][7]  ( .D(\row2_buffer[202][7] ), .CK(clk), .Q(
        \row2_buffer[201][7] ) );
  DFFQXL \row2_buffer_reg[200][7]  ( .D(\row2_buffer[201][7] ), .CK(clk), .Q(
        \row2_buffer[200][7] ) );
  DFFQXL \row2_buffer_reg[199][7]  ( .D(\row2_buffer[200][7] ), .CK(clk), .Q(
        \row2_buffer[199][7] ) );
  DFFQXL \row2_buffer_reg[198][7]  ( .D(\row2_buffer[199][7] ), .CK(clk), .Q(
        \row2_buffer[198][7] ) );
  DFFQXL \row2_buffer_reg[197][7]  ( .D(\row2_buffer[198][7] ), .CK(clk), .Q(
        \row2_buffer[197][7] ) );
  DFFQXL \row2_buffer_reg[196][7]  ( .D(\row2_buffer[197][7] ), .CK(clk), .Q(
        \row2_buffer[196][7] ) );
  DFFQXL \row2_buffer_reg[195][7]  ( .D(\row2_buffer[196][7] ), .CK(clk), .Q(
        \row2_buffer[195][7] ) );
  DFFQXL \row2_buffer_reg[194][7]  ( .D(\row2_buffer[195][7] ), .CK(clk), .Q(
        \row2_buffer[194][7] ) );
  DFFQXL \row2_buffer_reg[193][7]  ( .D(\row2_buffer[194][7] ), .CK(clk), .Q(
        \row2_buffer[193][7] ) );
  DFFQXL \row2_buffer_reg[192][7]  ( .D(\row2_buffer[193][7] ), .CK(clk), .Q(
        \row2_buffer[192][7] ) );
  DFFQXL \row2_buffer_reg[191][7]  ( .D(\row2_buffer[192][7] ), .CK(clk), .Q(
        \row2_buffer[191][7] ) );
  DFFQXL \row2_buffer_reg[190][7]  ( .D(\row2_buffer[191][7] ), .CK(clk), .Q(
        \row2_buffer[190][7] ) );
  DFFQXL \row2_buffer_reg[189][7]  ( .D(\row2_buffer[190][7] ), .CK(clk), .Q(
        \row2_buffer[189][7] ) );
  DFFQXL \row2_buffer_reg[188][7]  ( .D(\row2_buffer[189][7] ), .CK(clk), .Q(
        \row2_buffer[188][7] ) );
  DFFQXL \row2_buffer_reg[187][7]  ( .D(\row2_buffer[188][7] ), .CK(clk), .Q(
        \row2_buffer[187][7] ) );
  DFFQXL \row2_buffer_reg[186][7]  ( .D(\row2_buffer[187][7] ), .CK(clk), .Q(
        \row2_buffer[186][7] ) );
  DFFQXL \row2_buffer_reg[185][7]  ( .D(\row2_buffer[186][7] ), .CK(clk), .Q(
        \row2_buffer[185][7] ) );
  DFFQXL \row2_buffer_reg[184][7]  ( .D(\row2_buffer[185][7] ), .CK(clk), .Q(
        \row2_buffer[184][7] ) );
  DFFQXL \row2_buffer_reg[183][7]  ( .D(\row2_buffer[184][7] ), .CK(clk), .Q(
        \row2_buffer[183][7] ) );
  DFFQXL \row2_buffer_reg[182][7]  ( .D(\row2_buffer[183][7] ), .CK(clk), .Q(
        \row2_buffer[182][7] ) );
  DFFQXL \row2_buffer_reg[181][7]  ( .D(\row2_buffer[182][7] ), .CK(clk), .Q(
        \row2_buffer[181][7] ) );
  DFFQXL \row2_buffer_reg[180][7]  ( .D(\row2_buffer[181][7] ), .CK(clk), .Q(
        \row2_buffer[180][7] ) );
  DFFQXL \row2_buffer_reg[179][7]  ( .D(\row2_buffer[180][7] ), .CK(clk), .Q(
        \row2_buffer[179][7] ) );
  DFFQXL \row2_buffer_reg[178][7]  ( .D(\row2_buffer[179][7] ), .CK(clk), .Q(
        \row2_buffer[178][7] ) );
  DFFQXL \row2_buffer_reg[177][7]  ( .D(\row2_buffer[178][7] ), .CK(clk), .Q(
        \row2_buffer[177][7] ) );
  DFFQXL \row2_buffer_reg[176][7]  ( .D(\row2_buffer[177][7] ), .CK(clk), .Q(
        \row2_buffer[176][7] ) );
  DFFQXL \row2_buffer_reg[175][7]  ( .D(\row2_buffer[176][7] ), .CK(clk), .Q(
        \row2_buffer[175][7] ) );
  DFFQXL \row2_buffer_reg[174][7]  ( .D(\row2_buffer[175][7] ), .CK(clk), .Q(
        \row2_buffer[174][7] ) );
  DFFQXL \row2_buffer_reg[173][7]  ( .D(\row2_buffer[174][7] ), .CK(clk), .Q(
        \row2_buffer[173][7] ) );
  DFFQXL \row2_buffer_reg[172][7]  ( .D(\row2_buffer[173][7] ), .CK(clk), .Q(
        \row2_buffer[172][7] ) );
  DFFQXL \row2_buffer_reg[171][7]  ( .D(\row2_buffer[172][7] ), .CK(clk), .Q(
        \row2_buffer[171][7] ) );
  DFFQXL \row2_buffer_reg[170][7]  ( .D(\row2_buffer[171][7] ), .CK(clk), .Q(
        \row2_buffer[170][7] ) );
  DFFQXL \row2_buffer_reg[169][7]  ( .D(\row2_buffer[170][7] ), .CK(clk), .Q(
        \row2_buffer[169][7] ) );
  DFFQXL \row2_buffer_reg[168][7]  ( .D(\row2_buffer[169][7] ), .CK(clk), .Q(
        \row2_buffer[168][7] ) );
  DFFQXL \row2_buffer_reg[167][7]  ( .D(\row2_buffer[168][7] ), .CK(clk), .Q(
        \row2_buffer[167][7] ) );
  DFFQXL \row2_buffer_reg[166][7]  ( .D(\row2_buffer[167][7] ), .CK(clk), .Q(
        \row2_buffer[166][7] ) );
  DFFQXL \row2_buffer_reg[165][7]  ( .D(\row2_buffer[166][7] ), .CK(clk), .Q(
        \row2_buffer[165][7] ) );
  DFFQXL \row2_buffer_reg[164][7]  ( .D(\row2_buffer[165][7] ), .CK(clk), .Q(
        \row2_buffer[164][7] ) );
  DFFQXL \row2_buffer_reg[163][7]  ( .D(\row2_buffer[164][7] ), .CK(clk), .Q(
        \row2_buffer[163][7] ) );
  DFFQXL \row2_buffer_reg[162][7]  ( .D(\row2_buffer[163][7] ), .CK(clk), .Q(
        \row2_buffer[162][7] ) );
  DFFQXL \row2_buffer_reg[161][7]  ( .D(\row2_buffer[162][7] ), .CK(clk), .Q(
        \row2_buffer[161][7] ) );
  DFFQXL \row2_buffer_reg[160][7]  ( .D(\row2_buffer[161][7] ), .CK(clk), .Q(
        \row2_buffer[160][7] ) );
  DFFQXL \row2_buffer_reg[159][7]  ( .D(\row2_buffer[160][7] ), .CK(clk), .Q(
        \row2_buffer[159][7] ) );
  DFFQXL \row2_buffer_reg[158][7]  ( .D(\row2_buffer[159][7] ), .CK(clk), .Q(
        \row2_buffer[158][7] ) );
  DFFQXL \row2_buffer_reg[157][7]  ( .D(\row2_buffer[158][7] ), .CK(clk), .Q(
        \row2_buffer[157][7] ) );
  DFFQXL \row2_buffer_reg[156][7]  ( .D(\row2_buffer[157][7] ), .CK(clk), .Q(
        \row2_buffer[156][7] ) );
  DFFQXL \row2_buffer_reg[155][7]  ( .D(\row2_buffer[156][7] ), .CK(clk), .Q(
        \row2_buffer[155][7] ) );
  DFFQXL \row2_buffer_reg[154][7]  ( .D(\row2_buffer[155][7] ), .CK(clk), .Q(
        \row2_buffer[154][7] ) );
  DFFQXL \row2_buffer_reg[153][7]  ( .D(\row2_buffer[154][7] ), .CK(clk), .Q(
        \row2_buffer[153][7] ) );
  DFFQXL \row2_buffer_reg[152][7]  ( .D(\row2_buffer[153][7] ), .CK(clk), .Q(
        \row2_buffer[152][7] ) );
  DFFQXL \row2_buffer_reg[151][7]  ( .D(\row2_buffer[152][7] ), .CK(clk), .Q(
        \row2_buffer[151][7] ) );
  DFFQXL \row2_buffer_reg[150][7]  ( .D(\row2_buffer[151][7] ), .CK(clk), .Q(
        \row2_buffer[150][7] ) );
  DFFQXL \row2_buffer_reg[149][7]  ( .D(\row2_buffer[150][7] ), .CK(clk), .Q(
        \row2_buffer[149][7] ) );
  DFFQXL \row2_buffer_reg[148][7]  ( .D(\row2_buffer[149][7] ), .CK(clk), .Q(
        \row2_buffer[148][7] ) );
  DFFQXL \row2_buffer_reg[147][7]  ( .D(\row2_buffer[148][7] ), .CK(clk), .Q(
        \row2_buffer[147][7] ) );
  DFFQXL \row2_buffer_reg[146][7]  ( .D(\row2_buffer[147][7] ), .CK(clk), .Q(
        \row2_buffer[146][7] ) );
  DFFQXL \row2_buffer_reg[145][7]  ( .D(\row2_buffer[146][7] ), .CK(clk), .Q(
        \row2_buffer[145][7] ) );
  DFFQXL \row2_buffer_reg[144][7]  ( .D(\row2_buffer[145][7] ), .CK(clk), .Q(
        \row2_buffer[144][7] ) );
  DFFQXL \row2_buffer_reg[143][7]  ( .D(\row2_buffer[144][7] ), .CK(clk), .Q(
        \row2_buffer[143][7] ) );
  DFFQXL \row2_buffer_reg[142][7]  ( .D(\row2_buffer[143][7] ), .CK(clk), .Q(
        \row2_buffer[142][7] ) );
  DFFQXL \row2_buffer_reg[141][7]  ( .D(\row2_buffer[142][7] ), .CK(clk), .Q(
        \row2_buffer[141][7] ) );
  DFFQXL \row2_buffer_reg[140][7]  ( .D(\row2_buffer[141][7] ), .CK(clk), .Q(
        \row2_buffer[140][7] ) );
  DFFQXL \row2_buffer_reg[139][7]  ( .D(\row2_buffer[140][7] ), .CK(clk), .Q(
        \row2_buffer[139][7] ) );
  DFFQXL \row2_buffer_reg[138][7]  ( .D(\row2_buffer[139][7] ), .CK(clk), .Q(
        \row2_buffer[138][7] ) );
  DFFQXL \row2_buffer_reg[137][7]  ( .D(\row2_buffer[138][7] ), .CK(clk), .Q(
        \row2_buffer[137][7] ) );
  DFFQXL \row2_buffer_reg[136][7]  ( .D(\row2_buffer[137][7] ), .CK(clk), .Q(
        \row2_buffer[136][7] ) );
  DFFQXL \row2_buffer_reg[135][7]  ( .D(\row2_buffer[136][7] ), .CK(clk), .Q(
        \row2_buffer[135][7] ) );
  DFFQXL \row2_buffer_reg[134][7]  ( .D(\row2_buffer[135][7] ), .CK(clk), .Q(
        \row2_buffer[134][7] ) );
  DFFQXL \row2_buffer_reg[133][7]  ( .D(\row2_buffer[134][7] ), .CK(clk), .Q(
        \row2_buffer[133][7] ) );
  DFFQXL \row2_buffer_reg[132][7]  ( .D(\row2_buffer[133][7] ), .CK(clk), .Q(
        \row2_buffer[132][7] ) );
  DFFQXL \row2_buffer_reg[131][7]  ( .D(\row2_buffer[132][7] ), .CK(clk), .Q(
        \row2_buffer[131][7] ) );
  DFFQXL \row2_buffer_reg[130][7]  ( .D(\row2_buffer[131][7] ), .CK(clk), .Q(
        \row2_buffer[130][7] ) );
  DFFQXL \row2_buffer_reg[129][7]  ( .D(\row2_buffer[130][7] ), .CK(clk), .Q(
        \row2_buffer[129][7] ) );
  DFFQXL \row2_buffer_reg[128][7]  ( .D(\row2_buffer[129][7] ), .CK(clk), .Q(
        \row2_buffer[128][7] ) );
  DFFQXL \row2_buffer_reg[127][7]  ( .D(\row2_buffer[128][7] ), .CK(clk), .Q(
        \row2_buffer[127][7] ) );
  DFFQXL \row2_buffer_reg[126][7]  ( .D(\row2_buffer[127][7] ), .CK(clk), .Q(
        \row2_buffer[126][7] ) );
  DFFQXL \row2_buffer_reg[125][7]  ( .D(\row2_buffer[126][7] ), .CK(clk), .Q(
        \row2_buffer[125][7] ) );
  DFFQXL \row2_buffer_reg[124][7]  ( .D(\row2_buffer[125][7] ), .CK(clk), .Q(
        \row2_buffer[124][7] ) );
  DFFQXL \row2_buffer_reg[123][7]  ( .D(\row2_buffer[124][7] ), .CK(clk), .Q(
        \row2_buffer[123][7] ) );
  DFFQXL \row2_buffer_reg[122][7]  ( .D(\row2_buffer[123][7] ), .CK(clk), .Q(
        \row2_buffer[122][7] ) );
  DFFQXL \row2_buffer_reg[121][7]  ( .D(\row2_buffer[122][7] ), .CK(clk), .Q(
        \row2_buffer[121][7] ) );
  DFFQXL \row2_buffer_reg[120][7]  ( .D(\row2_buffer[121][7] ), .CK(clk), .Q(
        \row2_buffer[120][7] ) );
  DFFQXL \row2_buffer_reg[119][7]  ( .D(\row2_buffer[120][7] ), .CK(clk), .Q(
        \row2_buffer[119][7] ) );
  DFFQXL \row2_buffer_reg[118][7]  ( .D(\row2_buffer[119][7] ), .CK(clk), .Q(
        \row2_buffer[118][7] ) );
  DFFQXL \row2_buffer_reg[117][7]  ( .D(\row2_buffer[118][7] ), .CK(clk), .Q(
        \row2_buffer[117][7] ) );
  DFFQXL \row2_buffer_reg[116][7]  ( .D(\row2_buffer[117][7] ), .CK(clk), .Q(
        \row2_buffer[116][7] ) );
  DFFQXL \row2_buffer_reg[115][7]  ( .D(\row2_buffer[116][7] ), .CK(clk), .Q(
        \row2_buffer[115][7] ) );
  DFFQXL \row2_buffer_reg[114][7]  ( .D(\row2_buffer[115][7] ), .CK(clk), .Q(
        \row2_buffer[114][7] ) );
  DFFQXL \row2_buffer_reg[113][7]  ( .D(\row2_buffer[114][7] ), .CK(clk), .Q(
        \row2_buffer[113][7] ) );
  DFFQXL \row2_buffer_reg[112][7]  ( .D(\row2_buffer[113][7] ), .CK(clk), .Q(
        \row2_buffer[112][7] ) );
  DFFQXL \row2_buffer_reg[111][7]  ( .D(\row2_buffer[112][7] ), .CK(clk), .Q(
        \row2_buffer[111][7] ) );
  DFFQXL \row2_buffer_reg[110][7]  ( .D(\row2_buffer[111][7] ), .CK(clk), .Q(
        \row2_buffer[110][7] ) );
  DFFQXL \row2_buffer_reg[109][7]  ( .D(\row2_buffer[110][7] ), .CK(clk), .Q(
        \row2_buffer[109][7] ) );
  DFFQXL \row2_buffer_reg[108][7]  ( .D(\row2_buffer[109][7] ), .CK(clk), .Q(
        \row2_buffer[108][7] ) );
  DFFQXL \row2_buffer_reg[107][7]  ( .D(\row2_buffer[108][7] ), .CK(clk), .Q(
        \row2_buffer[107][7] ) );
  DFFQXL \row2_buffer_reg[106][7]  ( .D(\row2_buffer[107][7] ), .CK(clk), .Q(
        \row2_buffer[106][7] ) );
  DFFQXL \row2_buffer_reg[105][7]  ( .D(\row2_buffer[106][7] ), .CK(clk), .Q(
        \row2_buffer[105][7] ) );
  DFFQXL \row2_buffer_reg[104][7]  ( .D(\row2_buffer[105][7] ), .CK(clk), .Q(
        \row2_buffer[104][7] ) );
  DFFQXL \row2_buffer_reg[103][7]  ( .D(\row2_buffer[104][7] ), .CK(clk), .Q(
        \row2_buffer[103][7] ) );
  DFFQXL \row2_buffer_reg[102][7]  ( .D(\row2_buffer[103][7] ), .CK(clk), .Q(
        \row2_buffer[102][7] ) );
  DFFQXL \row2_buffer_reg[101][7]  ( .D(\row2_buffer[102][7] ), .CK(clk), .Q(
        \row2_buffer[101][7] ) );
  DFFQXL \row2_buffer_reg[100][7]  ( .D(\row2_buffer[101][7] ), .CK(clk), .Q(
        \row2_buffer[100][7] ) );
  DFFQXL \row2_buffer_reg[99][7]  ( .D(\row2_buffer[100][7] ), .CK(clk), .Q(
        \row2_buffer[99][7] ) );
  DFFQXL \row2_buffer_reg[98][7]  ( .D(\row2_buffer[99][7] ), .CK(clk), .Q(
        \row2_buffer[98][7] ) );
  DFFQXL \row2_buffer_reg[97][7]  ( .D(\row2_buffer[98][7] ), .CK(clk), .Q(
        \row2_buffer[97][7] ) );
  DFFQXL \row2_buffer_reg[96][7]  ( .D(\row2_buffer[97][7] ), .CK(clk), .Q(
        \row2_buffer[96][7] ) );
  DFFQXL \row2_buffer_reg[95][7]  ( .D(\row2_buffer[96][7] ), .CK(clk), .Q(
        \row2_buffer[95][7] ) );
  DFFQXL \row2_buffer_reg[94][7]  ( .D(\row2_buffer[95][7] ), .CK(clk), .Q(
        \row2_buffer[94][7] ) );
  DFFQXL \row2_buffer_reg[93][7]  ( .D(\row2_buffer[94][7] ), .CK(clk), .Q(
        \row2_buffer[93][7] ) );
  DFFQXL \row2_buffer_reg[92][7]  ( .D(\row2_buffer[93][7] ), .CK(clk), .Q(
        \row2_buffer[92][7] ) );
  DFFQXL \row2_buffer_reg[91][7]  ( .D(\row2_buffer[92][7] ), .CK(clk), .Q(
        \row2_buffer[91][7] ) );
  DFFQXL \row2_buffer_reg[90][7]  ( .D(\row2_buffer[91][7] ), .CK(clk), .Q(
        \row2_buffer[90][7] ) );
  DFFQXL \row2_buffer_reg[89][7]  ( .D(\row2_buffer[90][7] ), .CK(clk), .Q(
        \row2_buffer[89][7] ) );
  DFFQXL \row2_buffer_reg[88][7]  ( .D(\row2_buffer[89][7] ), .CK(clk), .Q(
        \row2_buffer[88][7] ) );
  DFFQXL \row2_buffer_reg[87][7]  ( .D(\row2_buffer[88][7] ), .CK(clk), .Q(
        \row2_buffer[87][7] ) );
  DFFQXL \row2_buffer_reg[86][7]  ( .D(\row2_buffer[87][7] ), .CK(clk), .Q(
        \row2_buffer[86][7] ) );
  DFFQXL \row2_buffer_reg[85][7]  ( .D(\row2_buffer[86][7] ), .CK(clk), .Q(
        \row2_buffer[85][7] ) );
  DFFQXL \row2_buffer_reg[84][7]  ( .D(\row2_buffer[85][7] ), .CK(clk), .Q(
        \row2_buffer[84][7] ) );
  DFFQXL \row2_buffer_reg[83][7]  ( .D(\row2_buffer[84][7] ), .CK(clk), .Q(
        \row2_buffer[83][7] ) );
  DFFQXL \row2_buffer_reg[82][7]  ( .D(\row2_buffer[83][7] ), .CK(clk), .Q(
        \row2_buffer[82][7] ) );
  DFFQXL \row2_buffer_reg[81][7]  ( .D(\row2_buffer[82][7] ), .CK(clk), .Q(
        \row2_buffer[81][7] ) );
  DFFQXL \row2_buffer_reg[80][7]  ( .D(\row2_buffer[81][7] ), .CK(clk), .Q(
        \row2_buffer[80][7] ) );
  DFFQXL \row2_buffer_reg[79][7]  ( .D(\row2_buffer[80][7] ), .CK(clk), .Q(
        \row2_buffer[79][7] ) );
  DFFQXL \row2_buffer_reg[78][7]  ( .D(\row2_buffer[79][7] ), .CK(clk), .Q(
        \row2_buffer[78][7] ) );
  DFFQXL \row2_buffer_reg[77][7]  ( .D(\row2_buffer[78][7] ), .CK(clk), .Q(
        \row2_buffer[77][7] ) );
  DFFQXL \row2_buffer_reg[76][7]  ( .D(\row2_buffer[77][7] ), .CK(clk), .Q(
        \row2_buffer[76][7] ) );
  DFFQXL \row2_buffer_reg[75][7]  ( .D(\row2_buffer[76][7] ), .CK(clk), .Q(
        \row2_buffer[75][7] ) );
  DFFQXL \row2_buffer_reg[74][7]  ( .D(\row2_buffer[75][7] ), .CK(clk), .Q(
        \row2_buffer[74][7] ) );
  DFFQXL \row2_buffer_reg[73][7]  ( .D(\row2_buffer[74][7] ), .CK(clk), .Q(
        \row2_buffer[73][7] ) );
  DFFQXL \row2_buffer_reg[72][7]  ( .D(\row2_buffer[73][7] ), .CK(clk), .Q(
        \row2_buffer[72][7] ) );
  DFFQXL \row2_buffer_reg[71][7]  ( .D(\row2_buffer[72][7] ), .CK(clk), .Q(
        \row2_buffer[71][7] ) );
  DFFQXL \row2_buffer_reg[70][7]  ( .D(\row2_buffer[71][7] ), .CK(clk), .Q(
        \row2_buffer[70][7] ) );
  DFFQXL \row2_buffer_reg[69][7]  ( .D(\row2_buffer[70][7] ), .CK(clk), .Q(
        \row2_buffer[69][7] ) );
  DFFQXL \row2_buffer_reg[68][7]  ( .D(\row2_buffer[69][7] ), .CK(clk), .Q(
        \row2_buffer[68][7] ) );
  DFFQXL \row2_buffer_reg[67][7]  ( .D(\row2_buffer[68][7] ), .CK(clk), .Q(
        \row2_buffer[67][7] ) );
  DFFQXL \row2_buffer_reg[66][7]  ( .D(\row2_buffer[67][7] ), .CK(clk), .Q(
        \row2_buffer[66][7] ) );
  DFFQXL \row2_buffer_reg[65][7]  ( .D(\row2_buffer[66][7] ), .CK(clk), .Q(
        \row2_buffer[65][7] ) );
  DFFQXL \row2_buffer_reg[64][7]  ( .D(\row2_buffer[65][7] ), .CK(clk), .Q(
        \row2_buffer[64][7] ) );
  DFFQXL \row2_buffer_reg[63][7]  ( .D(\row2_buffer[64][7] ), .CK(clk), .Q(
        \row2_buffer[63][7] ) );
  DFFQXL \row2_buffer_reg[62][7]  ( .D(\row2_buffer[63][7] ), .CK(clk), .Q(
        \row2_buffer[62][7] ) );
  DFFQXL \row2_buffer_reg[61][7]  ( .D(\row2_buffer[62][7] ), .CK(clk), .Q(
        \row2_buffer[61][7] ) );
  DFFQXL \row2_buffer_reg[60][7]  ( .D(\row2_buffer[61][7] ), .CK(clk), .Q(
        \row2_buffer[60][7] ) );
  DFFQXL \row2_buffer_reg[59][7]  ( .D(\row2_buffer[60][7] ), .CK(clk), .Q(
        \row2_buffer[59][7] ) );
  DFFQXL \row2_buffer_reg[58][7]  ( .D(\row2_buffer[59][7] ), .CK(clk), .Q(
        \row2_buffer[58][7] ) );
  DFFQXL \row2_buffer_reg[57][7]  ( .D(\row2_buffer[58][7] ), .CK(clk), .Q(
        \row2_buffer[57][7] ) );
  DFFQXL \row2_buffer_reg[56][7]  ( .D(\row2_buffer[57][7] ), .CK(clk), .Q(
        \row2_buffer[56][7] ) );
  DFFQXL \row2_buffer_reg[55][7]  ( .D(\row2_buffer[56][7] ), .CK(clk), .Q(
        \row2_buffer[55][7] ) );
  DFFQXL \row2_buffer_reg[54][7]  ( .D(\row2_buffer[55][7] ), .CK(clk), .Q(
        \row2_buffer[54][7] ) );
  DFFQXL \row2_buffer_reg[53][7]  ( .D(\row2_buffer[54][7] ), .CK(clk), .Q(
        \row2_buffer[53][7] ) );
  DFFQXL \row2_buffer_reg[52][7]  ( .D(\row2_buffer[53][7] ), .CK(clk), .Q(
        \row2_buffer[52][7] ) );
  DFFQXL \row2_buffer_reg[51][7]  ( .D(\row2_buffer[52][7] ), .CK(clk), .Q(
        \row2_buffer[51][7] ) );
  DFFQXL \row2_buffer_reg[50][7]  ( .D(\row2_buffer[51][7] ), .CK(clk), .Q(
        \row2_buffer[50][7] ) );
  DFFQXL \row2_buffer_reg[49][7]  ( .D(\row2_buffer[50][7] ), .CK(clk), .Q(
        \row2_buffer[49][7] ) );
  DFFQXL \row2_buffer_reg[48][7]  ( .D(\row2_buffer[49][7] ), .CK(clk), .Q(
        \row2_buffer[48][7] ) );
  DFFQXL \row2_buffer_reg[47][7]  ( .D(\row2_buffer[48][7] ), .CK(clk), .Q(
        \row2_buffer[47][7] ) );
  DFFQXL \row2_buffer_reg[46][7]  ( .D(\row2_buffer[47][7] ), .CK(clk), .Q(
        \row2_buffer[46][7] ) );
  DFFQXL \row2_buffer_reg[45][7]  ( .D(\row2_buffer[46][7] ), .CK(clk), .Q(
        \row2_buffer[45][7] ) );
  DFFQXL \row2_buffer_reg[44][7]  ( .D(\row2_buffer[45][7] ), .CK(clk), .Q(
        \row2_buffer[44][7] ) );
  DFFQXL \row2_buffer_reg[43][7]  ( .D(\row2_buffer[44][7] ), .CK(clk), .Q(
        \row2_buffer[43][7] ) );
  DFFQXL \row2_buffer_reg[42][7]  ( .D(\row2_buffer[43][7] ), .CK(clk), .Q(
        \row2_buffer[42][7] ) );
  DFFQXL \row2_buffer_reg[41][7]  ( .D(\row2_buffer[42][7] ), .CK(clk), .Q(
        \row2_buffer[41][7] ) );
  DFFQXL \row2_buffer_reg[40][7]  ( .D(\row2_buffer[41][7] ), .CK(clk), .Q(
        \row2_buffer[40][7] ) );
  DFFQXL \row2_buffer_reg[39][7]  ( .D(\row2_buffer[40][7] ), .CK(clk), .Q(
        \row2_buffer[39][7] ) );
  DFFQXL \row2_buffer_reg[38][7]  ( .D(\row2_buffer[39][7] ), .CK(clk), .Q(
        \row2_buffer[38][7] ) );
  DFFQXL \row2_buffer_reg[37][7]  ( .D(\row2_buffer[38][7] ), .CK(clk), .Q(
        \row2_buffer[37][7] ) );
  DFFQXL \row2_buffer_reg[36][7]  ( .D(\row2_buffer[37][7] ), .CK(clk), .Q(
        \row2_buffer[36][7] ) );
  DFFQXL \row2_buffer_reg[35][7]  ( .D(\row2_buffer[36][7] ), .CK(clk), .Q(
        \row2_buffer[35][7] ) );
  DFFQXL \row2_buffer_reg[34][7]  ( .D(\row2_buffer[35][7] ), .CK(clk), .Q(
        \row2_buffer[34][7] ) );
  DFFQXL \row2_buffer_reg[33][7]  ( .D(\row2_buffer[34][7] ), .CK(clk), .Q(
        \row2_buffer[33][7] ) );
  DFFQXL \row2_buffer_reg[32][7]  ( .D(\row2_buffer[33][7] ), .CK(clk), .Q(
        \row2_buffer[32][7] ) );
  DFFQXL \row2_buffer_reg[31][7]  ( .D(\row2_buffer[32][7] ), .CK(clk), .Q(
        \row2_buffer[31][7] ) );
  DFFQXL \row2_buffer_reg[30][7]  ( .D(\row2_buffer[31][7] ), .CK(clk), .Q(
        \row2_buffer[30][7] ) );
  DFFQXL \row2_buffer_reg[29][7]  ( .D(\row2_buffer[30][7] ), .CK(clk), .Q(
        \row2_buffer[29][7] ) );
  DFFQXL \row2_buffer_reg[28][7]  ( .D(\row2_buffer[29][7] ), .CK(clk), .Q(
        \row2_buffer[28][7] ) );
  DFFQXL \row2_buffer_reg[27][7]  ( .D(\row2_buffer[28][7] ), .CK(clk), .Q(
        \row2_buffer[27][7] ) );
  DFFQXL \row2_buffer_reg[26][7]  ( .D(\row2_buffer[27][7] ), .CK(clk), .Q(
        \row2_buffer[26][7] ) );
  DFFQXL \row2_buffer_reg[25][7]  ( .D(\row2_buffer[26][7] ), .CK(clk), .Q(
        \row2_buffer[25][7] ) );
  DFFQXL \row2_buffer_reg[24][7]  ( .D(\row2_buffer[25][7] ), .CK(clk), .Q(
        \row2_buffer[24][7] ) );
  DFFQXL \row2_buffer_reg[23][7]  ( .D(\row2_buffer[24][7] ), .CK(clk), .Q(
        \row2_buffer[23][7] ) );
  DFFQXL \row2_buffer_reg[22][7]  ( .D(\row2_buffer[23][7] ), .CK(clk), .Q(
        \row2_buffer[22][7] ) );
  DFFQXL \row2_buffer_reg[21][7]  ( .D(\row2_buffer[22][7] ), .CK(clk), .Q(
        \row2_buffer[21][7] ) );
  DFFQXL \row2_buffer_reg[20][7]  ( .D(\row2_buffer[21][7] ), .CK(clk), .Q(
        \row2_buffer[20][7] ) );
  DFFQXL \row2_buffer_reg[19][7]  ( .D(\row2_buffer[20][7] ), .CK(clk), .Q(
        \row2_buffer[19][7] ) );
  DFFQXL \row2_buffer_reg[18][7]  ( .D(\row2_buffer[19][7] ), .CK(clk), .Q(
        \row2_buffer[18][7] ) );
  DFFQXL \row2_buffer_reg[17][7]  ( .D(\row2_buffer[18][7] ), .CK(clk), .Q(
        \row2_buffer[17][7] ) );
  DFFQXL \row2_buffer_reg[16][7]  ( .D(\row2_buffer[17][7] ), .CK(clk), .Q(
        \row2_buffer[16][7] ) );
  DFFQXL \row2_buffer_reg[15][7]  ( .D(\row2_buffer[16][7] ), .CK(clk), .Q(
        \row2_buffer[15][7] ) );
  DFFQXL \row2_buffer_reg[14][7]  ( .D(\row2_buffer[15][7] ), .CK(clk), .Q(
        \row2_buffer[14][7] ) );
  DFFQXL \row2_buffer_reg[13][7]  ( .D(\row2_buffer[14][7] ), .CK(clk), .Q(
        \row2_buffer[13][7] ) );
  DFFQXL \row2_buffer_reg[12][7]  ( .D(\row2_buffer[13][7] ), .CK(clk), .Q(
        \row2_buffer[12][7] ) );
  DFFQXL \row2_buffer_reg[11][7]  ( .D(\row2_buffer[12][7] ), .CK(clk), .Q(
        \row2_buffer[11][7] ) );
  DFFQXL \row2_buffer_reg[10][7]  ( .D(\row2_buffer[11][7] ), .CK(clk), .Q(
        \row2_buffer[10][7] ) );
  DFFQXL \row2_buffer_reg[9][7]  ( .D(\row2_buffer[10][7] ), .CK(clk), .Q(
        \row2_buffer[9][7] ) );
  DFFQXL \row2_buffer_reg[8][7]  ( .D(\row2_buffer[9][7] ), .CK(clk), .Q(
        \row2_buffer[8][7] ) );
  DFFQXL \row2_buffer_reg[7][7]  ( .D(\row2_buffer[8][7] ), .CK(clk), .Q(
        \row2_buffer[7][7] ) );
  DFFQXL \row2_buffer_reg[6][7]  ( .D(\row2_buffer[7][7] ), .CK(clk), .Q(
        \row2_buffer[6][7] ) );
  DFFQXL \row2_buffer_reg[5][7]  ( .D(\row2_buffer[6][7] ), .CK(clk), .Q(
        \row2_buffer[5][7] ) );
  DFFQXL \row2_buffer_reg[4][7]  ( .D(\row2_buffer[5][7] ), .CK(clk), .Q(
        \row2_buffer[4][7] ) );
  DFFQXL \row2_buffer_reg[3][7]  ( .D(\row2_buffer[4][7] ), .CK(clk), .Q(
        \row2_buffer[3][7] ) );
  DFFQXL \row1_buffer_reg[225][7]  ( .D(\row2_buffer[0][7] ), .CK(clk), .Q(
        \row1_buffer[225][7] ) );
  DFFQXL \row1_buffer_reg[224][7]  ( .D(\row1_buffer[225][7] ), .CK(clk), .Q(
        \row1_buffer[224][7] ) );
  DFFQXL \row1_buffer_reg[223][7]  ( .D(\row1_buffer[224][7] ), .CK(clk), .Q(
        \row1_buffer[223][7] ) );
  DFFQXL \row1_buffer_reg[222][7]  ( .D(\row1_buffer[223][7] ), .CK(clk), .Q(
        \row1_buffer[222][7] ) );
  DFFQXL \row1_buffer_reg[221][7]  ( .D(\row1_buffer[222][7] ), .CK(clk), .Q(
        \row1_buffer[221][7] ) );
  DFFQXL \row1_buffer_reg[220][7]  ( .D(\row1_buffer[221][7] ), .CK(clk), .Q(
        \row1_buffer[220][7] ) );
  DFFQXL \row1_buffer_reg[219][7]  ( .D(\row1_buffer[220][7] ), .CK(clk), .Q(
        \row1_buffer[219][7] ) );
  DFFQXL \row1_buffer_reg[218][7]  ( .D(\row1_buffer[219][7] ), .CK(clk), .Q(
        \row1_buffer[218][7] ) );
  DFFQXL \row1_buffer_reg[217][7]  ( .D(\row1_buffer[218][7] ), .CK(clk), .Q(
        \row1_buffer[217][7] ) );
  DFFQXL \row1_buffer_reg[216][7]  ( .D(\row1_buffer[217][7] ), .CK(clk), .Q(
        \row1_buffer[216][7] ) );
  DFFQXL \row1_buffer_reg[215][7]  ( .D(\row1_buffer[216][7] ), .CK(clk), .Q(
        \row1_buffer[215][7] ) );
  DFFQXL \row1_buffer_reg[214][7]  ( .D(\row1_buffer[215][7] ), .CK(clk), .Q(
        \row1_buffer[214][7] ) );
  DFFQXL \row1_buffer_reg[213][7]  ( .D(\row1_buffer[214][7] ), .CK(clk), .Q(
        \row1_buffer[213][7] ) );
  DFFQXL \row1_buffer_reg[212][7]  ( .D(\row1_buffer[213][7] ), .CK(clk), .Q(
        \row1_buffer[212][7] ) );
  DFFQXL \row1_buffer_reg[211][7]  ( .D(\row1_buffer[212][7] ), .CK(clk), .Q(
        \row1_buffer[211][7] ) );
  DFFQXL \row1_buffer_reg[210][7]  ( .D(\row1_buffer[211][7] ), .CK(clk), .Q(
        \row1_buffer[210][7] ) );
  DFFQXL \row1_buffer_reg[209][7]  ( .D(\row1_buffer[210][7] ), .CK(clk), .Q(
        \row1_buffer[209][7] ) );
  DFFQXL \row1_buffer_reg[208][7]  ( .D(\row1_buffer[209][7] ), .CK(clk), .Q(
        \row1_buffer[208][7] ) );
  DFFQXL \row1_buffer_reg[207][7]  ( .D(\row1_buffer[208][7] ), .CK(clk), .Q(
        \row1_buffer[207][7] ) );
  DFFQXL \row1_buffer_reg[206][7]  ( .D(\row1_buffer[207][7] ), .CK(clk), .Q(
        \row1_buffer[206][7] ) );
  DFFQXL \row1_buffer_reg[205][7]  ( .D(\row1_buffer[206][7] ), .CK(clk), .Q(
        \row1_buffer[205][7] ) );
  DFFQXL \row1_buffer_reg[204][7]  ( .D(\row1_buffer[205][7] ), .CK(clk), .Q(
        \row1_buffer[204][7] ) );
  DFFQXL \row1_buffer_reg[203][7]  ( .D(\row1_buffer[204][7] ), .CK(clk), .Q(
        \row1_buffer[203][7] ) );
  DFFQXL \row1_buffer_reg[202][7]  ( .D(\row1_buffer[203][7] ), .CK(clk), .Q(
        \row1_buffer[202][7] ) );
  DFFQXL \row1_buffer_reg[201][7]  ( .D(\row1_buffer[202][7] ), .CK(clk), .Q(
        \row1_buffer[201][7] ) );
  DFFQXL \row1_buffer_reg[200][7]  ( .D(\row1_buffer[201][7] ), .CK(clk), .Q(
        \row1_buffer[200][7] ) );
  DFFQXL \row1_buffer_reg[199][7]  ( .D(\row1_buffer[200][7] ), .CK(clk), .Q(
        \row1_buffer[199][7] ) );
  DFFQXL \row1_buffer_reg[198][7]  ( .D(\row1_buffer[199][7] ), .CK(clk), .Q(
        \row1_buffer[198][7] ) );
  DFFQXL \row1_buffer_reg[197][7]  ( .D(\row1_buffer[198][7] ), .CK(clk), .Q(
        \row1_buffer[197][7] ) );
  DFFQXL \row1_buffer_reg[196][7]  ( .D(\row1_buffer[197][7] ), .CK(clk), .Q(
        \row1_buffer[196][7] ) );
  DFFQXL \row1_buffer_reg[195][7]  ( .D(\row1_buffer[196][7] ), .CK(clk), .Q(
        \row1_buffer[195][7] ) );
  DFFQXL \row1_buffer_reg[194][7]  ( .D(\row1_buffer[195][7] ), .CK(clk), .Q(
        \row1_buffer[194][7] ) );
  DFFQXL \row1_buffer_reg[193][7]  ( .D(\row1_buffer[194][7] ), .CK(clk), .Q(
        \row1_buffer[193][7] ) );
  DFFQXL \row1_buffer_reg[192][7]  ( .D(\row1_buffer[193][7] ), .CK(clk), .Q(
        \row1_buffer[192][7] ) );
  DFFQXL \row1_buffer_reg[191][7]  ( .D(\row1_buffer[192][7] ), .CK(clk), .Q(
        \row1_buffer[191][7] ) );
  DFFQXL \row1_buffer_reg[190][7]  ( .D(\row1_buffer[191][7] ), .CK(clk), .Q(
        \row1_buffer[190][7] ) );
  DFFQXL \row1_buffer_reg[189][7]  ( .D(\row1_buffer[190][7] ), .CK(clk), .Q(
        \row1_buffer[189][7] ) );
  DFFQXL \row1_buffer_reg[188][7]  ( .D(\row1_buffer[189][7] ), .CK(clk), .Q(
        \row1_buffer[188][7] ) );
  DFFQXL \row1_buffer_reg[187][7]  ( .D(\row1_buffer[188][7] ), .CK(clk), .Q(
        \row1_buffer[187][7] ) );
  DFFQXL \row1_buffer_reg[186][7]  ( .D(\row1_buffer[187][7] ), .CK(clk), .Q(
        \row1_buffer[186][7] ) );
  DFFQXL \row1_buffer_reg[185][7]  ( .D(\row1_buffer[186][7] ), .CK(clk), .Q(
        \row1_buffer[185][7] ) );
  DFFQXL \row1_buffer_reg[184][7]  ( .D(\row1_buffer[185][7] ), .CK(clk), .Q(
        \row1_buffer[184][7] ) );
  DFFQXL \row1_buffer_reg[183][7]  ( .D(\row1_buffer[184][7] ), .CK(clk), .Q(
        \row1_buffer[183][7] ) );
  DFFQXL \row1_buffer_reg[182][7]  ( .D(\row1_buffer[183][7] ), .CK(clk), .Q(
        \row1_buffer[182][7] ) );
  DFFQXL \row1_buffer_reg[181][7]  ( .D(\row1_buffer[182][7] ), .CK(clk), .Q(
        \row1_buffer[181][7] ) );
  DFFQXL \row1_buffer_reg[180][7]  ( .D(\row1_buffer[181][7] ), .CK(clk), .Q(
        \row1_buffer[180][7] ) );
  DFFQXL \row1_buffer_reg[179][7]  ( .D(\row1_buffer[180][7] ), .CK(clk), .Q(
        \row1_buffer[179][7] ) );
  DFFQXL \row1_buffer_reg[178][7]  ( .D(\row1_buffer[179][7] ), .CK(clk), .Q(
        \row1_buffer[178][7] ) );
  DFFQXL \row1_buffer_reg[177][7]  ( .D(\row1_buffer[178][7] ), .CK(clk), .Q(
        \row1_buffer[177][7] ) );
  DFFQXL \row1_buffer_reg[176][7]  ( .D(\row1_buffer[177][7] ), .CK(clk), .Q(
        \row1_buffer[176][7] ) );
  DFFQXL \row1_buffer_reg[175][7]  ( .D(\row1_buffer[176][7] ), .CK(clk), .Q(
        \row1_buffer[175][7] ) );
  DFFQXL \row1_buffer_reg[174][7]  ( .D(\row1_buffer[175][7] ), .CK(clk), .Q(
        \row1_buffer[174][7] ) );
  DFFQXL \row1_buffer_reg[173][7]  ( .D(\row1_buffer[174][7] ), .CK(clk), .Q(
        \row1_buffer[173][7] ) );
  DFFQXL \row1_buffer_reg[172][7]  ( .D(\row1_buffer[173][7] ), .CK(clk), .Q(
        \row1_buffer[172][7] ) );
  DFFQXL \row1_buffer_reg[171][7]  ( .D(\row1_buffer[172][7] ), .CK(clk), .Q(
        \row1_buffer[171][7] ) );
  DFFQXL \row1_buffer_reg[170][7]  ( .D(\row1_buffer[171][7] ), .CK(clk), .Q(
        \row1_buffer[170][7] ) );
  DFFQXL \row1_buffer_reg[169][7]  ( .D(\row1_buffer[170][7] ), .CK(clk), .Q(
        \row1_buffer[169][7] ) );
  DFFQXL \row1_buffer_reg[168][7]  ( .D(\row1_buffer[169][7] ), .CK(clk), .Q(
        \row1_buffer[168][7] ) );
  DFFQXL \row1_buffer_reg[167][7]  ( .D(\row1_buffer[168][7] ), .CK(clk), .Q(
        \row1_buffer[167][7] ) );
  DFFQXL \row1_buffer_reg[166][7]  ( .D(\row1_buffer[167][7] ), .CK(clk), .Q(
        \row1_buffer[166][7] ) );
  DFFQXL \row1_buffer_reg[165][7]  ( .D(\row1_buffer[166][7] ), .CK(clk), .Q(
        \row1_buffer[165][7] ) );
  DFFQXL \row1_buffer_reg[164][7]  ( .D(\row1_buffer[165][7] ), .CK(clk), .Q(
        \row1_buffer[164][7] ) );
  DFFQXL \row1_buffer_reg[163][7]  ( .D(\row1_buffer[164][7] ), .CK(clk), .Q(
        \row1_buffer[163][7] ) );
  DFFQXL \row1_buffer_reg[162][7]  ( .D(\row1_buffer[163][7] ), .CK(clk), .Q(
        \row1_buffer[162][7] ) );
  DFFQXL \row1_buffer_reg[161][7]  ( .D(\row1_buffer[162][7] ), .CK(clk), .Q(
        \row1_buffer[161][7] ) );
  DFFQXL \row1_buffer_reg[160][7]  ( .D(\row1_buffer[161][7] ), .CK(clk), .Q(
        \row1_buffer[160][7] ) );
  DFFQXL \row1_buffer_reg[159][7]  ( .D(\row1_buffer[160][7] ), .CK(clk), .Q(
        \row1_buffer[159][7] ) );
  DFFQXL \row1_buffer_reg[158][7]  ( .D(\row1_buffer[159][7] ), .CK(clk), .Q(
        \row1_buffer[158][7] ) );
  DFFQXL \row1_buffer_reg[157][7]  ( .D(\row1_buffer[158][7] ), .CK(clk), .Q(
        \row1_buffer[157][7] ) );
  DFFQXL \row1_buffer_reg[156][7]  ( .D(\row1_buffer[157][7] ), .CK(clk), .Q(
        \row1_buffer[156][7] ) );
  DFFQXL \row1_buffer_reg[155][7]  ( .D(\row1_buffer[156][7] ), .CK(clk), .Q(
        \row1_buffer[155][7] ) );
  DFFQXL \row1_buffer_reg[154][7]  ( .D(\row1_buffer[155][7] ), .CK(clk), .Q(
        \row1_buffer[154][7] ) );
  DFFQXL \row1_buffer_reg[153][7]  ( .D(\row1_buffer[154][7] ), .CK(clk), .Q(
        \row1_buffer[153][7] ) );
  DFFQXL \row1_buffer_reg[152][7]  ( .D(\row1_buffer[153][7] ), .CK(clk), .Q(
        \row1_buffer[152][7] ) );
  DFFQXL \row1_buffer_reg[151][7]  ( .D(\row1_buffer[152][7] ), .CK(clk), .Q(
        \row1_buffer[151][7] ) );
  DFFQXL \row1_buffer_reg[150][7]  ( .D(\row1_buffer[151][7] ), .CK(clk), .Q(
        \row1_buffer[150][7] ) );
  DFFQXL \row1_buffer_reg[149][7]  ( .D(\row1_buffer[150][7] ), .CK(clk), .Q(
        \row1_buffer[149][7] ) );
  DFFQXL \row1_buffer_reg[148][7]  ( .D(\row1_buffer[149][7] ), .CK(clk), .Q(
        \row1_buffer[148][7] ) );
  DFFQXL \row1_buffer_reg[147][7]  ( .D(\row1_buffer[148][7] ), .CK(clk), .Q(
        \row1_buffer[147][7] ) );
  DFFQXL \row1_buffer_reg[146][7]  ( .D(\row1_buffer[147][7] ), .CK(clk), .Q(
        \row1_buffer[146][7] ) );
  DFFQXL \row1_buffer_reg[145][7]  ( .D(\row1_buffer[146][7] ), .CK(clk), .Q(
        \row1_buffer[145][7] ) );
  DFFQXL \row1_buffer_reg[144][7]  ( .D(\row1_buffer[145][7] ), .CK(clk), .Q(
        \row1_buffer[144][7] ) );
  DFFQXL \row1_buffer_reg[143][7]  ( .D(\row1_buffer[144][7] ), .CK(clk), .Q(
        \row1_buffer[143][7] ) );
  DFFQXL \row1_buffer_reg[142][7]  ( .D(\row1_buffer[143][7] ), .CK(clk), .Q(
        \row1_buffer[142][7] ) );
  DFFQXL \row1_buffer_reg[141][7]  ( .D(\row1_buffer[142][7] ), .CK(clk), .Q(
        \row1_buffer[141][7] ) );
  DFFQXL \row1_buffer_reg[140][7]  ( .D(\row1_buffer[141][7] ), .CK(clk), .Q(
        \row1_buffer[140][7] ) );
  DFFQXL \row1_buffer_reg[139][7]  ( .D(\row1_buffer[140][7] ), .CK(clk), .Q(
        \row1_buffer[139][7] ) );
  DFFQXL \row1_buffer_reg[138][7]  ( .D(\row1_buffer[139][7] ), .CK(clk), .Q(
        \row1_buffer[138][7] ) );
  DFFQXL \row1_buffer_reg[137][7]  ( .D(\row1_buffer[138][7] ), .CK(clk), .Q(
        \row1_buffer[137][7] ) );
  DFFQXL \row1_buffer_reg[136][7]  ( .D(\row1_buffer[137][7] ), .CK(clk), .Q(
        \row1_buffer[136][7] ) );
  DFFQXL \row1_buffer_reg[135][7]  ( .D(\row1_buffer[136][7] ), .CK(clk), .Q(
        \row1_buffer[135][7] ) );
  DFFQXL \row1_buffer_reg[134][7]  ( .D(\row1_buffer[135][7] ), .CK(clk), .Q(
        \row1_buffer[134][7] ) );
  DFFQXL \row1_buffer_reg[133][7]  ( .D(\row1_buffer[134][7] ), .CK(clk), .Q(
        \row1_buffer[133][7] ) );
  DFFQXL \row1_buffer_reg[132][7]  ( .D(\row1_buffer[133][7] ), .CK(clk), .Q(
        \row1_buffer[132][7] ) );
  DFFQXL \row1_buffer_reg[131][7]  ( .D(\row1_buffer[132][7] ), .CK(clk), .Q(
        \row1_buffer[131][7] ) );
  DFFQXL \row1_buffer_reg[130][7]  ( .D(\row1_buffer[131][7] ), .CK(clk), .Q(
        \row1_buffer[130][7] ) );
  DFFQXL \row1_buffer_reg[129][7]  ( .D(\row1_buffer[130][7] ), .CK(clk), .Q(
        \row1_buffer[129][7] ) );
  DFFQXL \row1_buffer_reg[128][7]  ( .D(\row1_buffer[129][7] ), .CK(clk), .Q(
        \row1_buffer[128][7] ) );
  DFFQXL \row1_buffer_reg[127][7]  ( .D(\row1_buffer[128][7] ), .CK(clk), .Q(
        \row1_buffer[127][7] ) );
  DFFQXL \row1_buffer_reg[126][7]  ( .D(\row1_buffer[127][7] ), .CK(clk), .Q(
        \row1_buffer[126][7] ) );
  DFFQXL \row1_buffer_reg[125][7]  ( .D(\row1_buffer[126][7] ), .CK(clk), .Q(
        \row1_buffer[125][7] ) );
  DFFQXL \row1_buffer_reg[124][7]  ( .D(\row1_buffer[125][7] ), .CK(clk), .Q(
        \row1_buffer[124][7] ) );
  DFFQXL \row1_buffer_reg[123][7]  ( .D(\row1_buffer[124][7] ), .CK(clk), .Q(
        \row1_buffer[123][7] ) );
  DFFQXL \row1_buffer_reg[122][7]  ( .D(\row1_buffer[123][7] ), .CK(clk), .Q(
        \row1_buffer[122][7] ) );
  DFFQXL \row1_buffer_reg[121][7]  ( .D(\row1_buffer[122][7] ), .CK(clk), .Q(
        \row1_buffer[121][7] ) );
  DFFQXL \row1_buffer_reg[120][7]  ( .D(\row1_buffer[121][7] ), .CK(clk), .Q(
        \row1_buffer[120][7] ) );
  DFFQXL \row1_buffer_reg[119][7]  ( .D(\row1_buffer[120][7] ), .CK(clk), .Q(
        \row1_buffer[119][7] ) );
  DFFQXL \row1_buffer_reg[118][7]  ( .D(\row1_buffer[119][7] ), .CK(clk), .Q(
        \row1_buffer[118][7] ) );
  DFFQXL \row1_buffer_reg[117][7]  ( .D(\row1_buffer[118][7] ), .CK(clk), .Q(
        \row1_buffer[117][7] ) );
  DFFQXL \row1_buffer_reg[116][7]  ( .D(\row1_buffer[117][7] ), .CK(clk), .Q(
        \row1_buffer[116][7] ) );
  DFFQXL \row1_buffer_reg[115][7]  ( .D(\row1_buffer[116][7] ), .CK(clk), .Q(
        \row1_buffer[115][7] ) );
  DFFQXL \row1_buffer_reg[114][7]  ( .D(\row1_buffer[115][7] ), .CK(clk), .Q(
        \row1_buffer[114][7] ) );
  DFFQXL \row1_buffer_reg[113][7]  ( .D(\row1_buffer[114][7] ), .CK(clk), .Q(
        \row1_buffer[113][7] ) );
  DFFQXL \row1_buffer_reg[112][7]  ( .D(\row1_buffer[113][7] ), .CK(clk), .Q(
        \row1_buffer[112][7] ) );
  DFFQXL \row1_buffer_reg[111][7]  ( .D(\row1_buffer[112][7] ), .CK(clk), .Q(
        \row1_buffer[111][7] ) );
  DFFQXL \row1_buffer_reg[110][7]  ( .D(\row1_buffer[111][7] ), .CK(clk), .Q(
        \row1_buffer[110][7] ) );
  DFFQXL \row1_buffer_reg[109][7]  ( .D(\row1_buffer[110][7] ), .CK(clk), .Q(
        \row1_buffer[109][7] ) );
  DFFQXL \row1_buffer_reg[108][7]  ( .D(\row1_buffer[109][7] ), .CK(clk), .Q(
        \row1_buffer[108][7] ) );
  DFFQXL \row1_buffer_reg[107][7]  ( .D(\row1_buffer[108][7] ), .CK(clk), .Q(
        \row1_buffer[107][7] ) );
  DFFQXL \row1_buffer_reg[106][7]  ( .D(\row1_buffer[107][7] ), .CK(clk), .Q(
        \row1_buffer[106][7] ) );
  DFFQXL \row1_buffer_reg[105][7]  ( .D(\row1_buffer[106][7] ), .CK(clk), .Q(
        \row1_buffer[105][7] ) );
  DFFQXL \row1_buffer_reg[104][7]  ( .D(\row1_buffer[105][7] ), .CK(clk), .Q(
        \row1_buffer[104][7] ) );
  DFFQXL \row1_buffer_reg[103][7]  ( .D(\row1_buffer[104][7] ), .CK(clk), .Q(
        \row1_buffer[103][7] ) );
  DFFQXL \row1_buffer_reg[102][7]  ( .D(\row1_buffer[103][7] ), .CK(clk), .Q(
        \row1_buffer[102][7] ) );
  DFFQXL \row1_buffer_reg[101][7]  ( .D(\row1_buffer[102][7] ), .CK(clk), .Q(
        \row1_buffer[101][7] ) );
  DFFQXL \row1_buffer_reg[100][7]  ( .D(\row1_buffer[101][7] ), .CK(clk), .Q(
        \row1_buffer[100][7] ) );
  DFFQXL \row1_buffer_reg[99][7]  ( .D(\row1_buffer[100][7] ), .CK(clk), .Q(
        \row1_buffer[99][7] ) );
  DFFQXL \row1_buffer_reg[98][7]  ( .D(\row1_buffer[99][7] ), .CK(clk), .Q(
        \row1_buffer[98][7] ) );
  DFFQXL \row1_buffer_reg[97][7]  ( .D(\row1_buffer[98][7] ), .CK(clk), .Q(
        \row1_buffer[97][7] ) );
  DFFQXL \row1_buffer_reg[96][7]  ( .D(\row1_buffer[97][7] ), .CK(clk), .Q(
        \row1_buffer[96][7] ) );
  DFFQXL \row1_buffer_reg[95][7]  ( .D(\row1_buffer[96][7] ), .CK(clk), .Q(
        \row1_buffer[95][7] ) );
  DFFQXL \row1_buffer_reg[94][7]  ( .D(\row1_buffer[95][7] ), .CK(clk), .Q(
        \row1_buffer[94][7] ) );
  DFFQXL \row1_buffer_reg[93][7]  ( .D(\row1_buffer[94][7] ), .CK(clk), .Q(
        \row1_buffer[93][7] ) );
  DFFQXL \row1_buffer_reg[92][7]  ( .D(\row1_buffer[93][7] ), .CK(clk), .Q(
        \row1_buffer[92][7] ) );
  DFFQXL \row1_buffer_reg[91][7]  ( .D(\row1_buffer[92][7] ), .CK(clk), .Q(
        \row1_buffer[91][7] ) );
  DFFQXL \row1_buffer_reg[90][7]  ( .D(\row1_buffer[91][7] ), .CK(clk), .Q(
        \row1_buffer[90][7] ) );
  DFFQXL \row1_buffer_reg[89][7]  ( .D(\row1_buffer[90][7] ), .CK(clk), .Q(
        \row1_buffer[89][7] ) );
  DFFQXL \row1_buffer_reg[88][7]  ( .D(\row1_buffer[89][7] ), .CK(clk), .Q(
        \row1_buffer[88][7] ) );
  DFFQXL \row1_buffer_reg[87][7]  ( .D(\row1_buffer[88][7] ), .CK(clk), .Q(
        \row1_buffer[87][7] ) );
  DFFQXL \row1_buffer_reg[86][7]  ( .D(\row1_buffer[87][7] ), .CK(clk), .Q(
        \row1_buffer[86][7] ) );
  DFFQXL \row1_buffer_reg[85][7]  ( .D(\row1_buffer[86][7] ), .CK(clk), .Q(
        \row1_buffer[85][7] ) );
  DFFQXL \row1_buffer_reg[84][7]  ( .D(\row1_buffer[85][7] ), .CK(clk), .Q(
        \row1_buffer[84][7] ) );
  DFFQXL \row1_buffer_reg[83][7]  ( .D(\row1_buffer[84][7] ), .CK(clk), .Q(
        \row1_buffer[83][7] ) );
  DFFQXL \row1_buffer_reg[82][7]  ( .D(\row1_buffer[83][7] ), .CK(clk), .Q(
        \row1_buffer[82][7] ) );
  DFFQXL \row1_buffer_reg[81][7]  ( .D(\row1_buffer[82][7] ), .CK(clk), .Q(
        \row1_buffer[81][7] ) );
  DFFQXL \row1_buffer_reg[80][7]  ( .D(\row1_buffer[81][7] ), .CK(clk), .Q(
        \row1_buffer[80][7] ) );
  DFFQXL \row1_buffer_reg[79][7]  ( .D(\row1_buffer[80][7] ), .CK(clk), .Q(
        \row1_buffer[79][7] ) );
  DFFQXL \row1_buffer_reg[78][7]  ( .D(\row1_buffer[79][7] ), .CK(clk), .Q(
        \row1_buffer[78][7] ) );
  DFFQXL \row1_buffer_reg[77][7]  ( .D(\row1_buffer[78][7] ), .CK(clk), .Q(
        \row1_buffer[77][7] ) );
  DFFQXL \row1_buffer_reg[76][7]  ( .D(\row1_buffer[77][7] ), .CK(clk), .Q(
        \row1_buffer[76][7] ) );
  DFFQXL \row1_buffer_reg[75][7]  ( .D(\row1_buffer[76][7] ), .CK(clk), .Q(
        \row1_buffer[75][7] ) );
  DFFQXL \row1_buffer_reg[74][7]  ( .D(\row1_buffer[75][7] ), .CK(clk), .Q(
        \row1_buffer[74][7] ) );
  DFFQXL \row1_buffer_reg[73][7]  ( .D(\row1_buffer[74][7] ), .CK(clk), .Q(
        \row1_buffer[73][7] ) );
  DFFQXL \row1_buffer_reg[72][7]  ( .D(\row1_buffer[73][7] ), .CK(clk), .Q(
        \row1_buffer[72][7] ) );
  DFFQXL \row1_buffer_reg[71][7]  ( .D(\row1_buffer[72][7] ), .CK(clk), .Q(
        \row1_buffer[71][7] ) );
  DFFQXL \row1_buffer_reg[70][7]  ( .D(\row1_buffer[71][7] ), .CK(clk), .Q(
        \row1_buffer[70][7] ) );
  DFFQXL \row1_buffer_reg[69][7]  ( .D(\row1_buffer[70][7] ), .CK(clk), .Q(
        \row1_buffer[69][7] ) );
  DFFQXL \row1_buffer_reg[68][7]  ( .D(\row1_buffer[69][7] ), .CK(clk), .Q(
        \row1_buffer[68][7] ) );
  DFFQXL \row1_buffer_reg[67][7]  ( .D(\row1_buffer[68][7] ), .CK(clk), .Q(
        \row1_buffer[67][7] ) );
  DFFQXL \row1_buffer_reg[66][7]  ( .D(\row1_buffer[67][7] ), .CK(clk), .Q(
        \row1_buffer[66][7] ) );
  DFFQXL \row1_buffer_reg[65][7]  ( .D(\row1_buffer[66][7] ), .CK(clk), .Q(
        \row1_buffer[65][7] ) );
  DFFQXL \row1_buffer_reg[64][7]  ( .D(\row1_buffer[65][7] ), .CK(clk), .Q(
        \row1_buffer[64][7] ) );
  DFFQXL \row1_buffer_reg[63][7]  ( .D(\row1_buffer[64][7] ), .CK(clk), .Q(
        \row1_buffer[63][7] ) );
  DFFQXL \row1_buffer_reg[62][7]  ( .D(\row1_buffer[63][7] ), .CK(clk), .Q(
        \row1_buffer[62][7] ) );
  DFFQXL \row1_buffer_reg[61][7]  ( .D(\row1_buffer[62][7] ), .CK(clk), .Q(
        \row1_buffer[61][7] ) );
  DFFQXL \row1_buffer_reg[60][7]  ( .D(\row1_buffer[61][7] ), .CK(clk), .Q(
        \row1_buffer[60][7] ) );
  DFFQXL \row1_buffer_reg[59][7]  ( .D(\row1_buffer[60][7] ), .CK(clk), .Q(
        \row1_buffer[59][7] ) );
  DFFQXL \row1_buffer_reg[58][7]  ( .D(\row1_buffer[59][7] ), .CK(clk), .Q(
        \row1_buffer[58][7] ) );
  DFFQXL \row1_buffer_reg[57][7]  ( .D(\row1_buffer[58][7] ), .CK(clk), .Q(
        \row1_buffer[57][7] ) );
  DFFQXL \row1_buffer_reg[56][7]  ( .D(\row1_buffer[57][7] ), .CK(clk), .Q(
        \row1_buffer[56][7] ) );
  DFFQXL \row1_buffer_reg[55][7]  ( .D(\row1_buffer[56][7] ), .CK(clk), .Q(
        \row1_buffer[55][7] ) );
  DFFQXL \row1_buffer_reg[54][7]  ( .D(\row1_buffer[55][7] ), .CK(clk), .Q(
        \row1_buffer[54][7] ) );
  DFFQXL \row1_buffer_reg[53][7]  ( .D(\row1_buffer[54][7] ), .CK(clk), .Q(
        \row1_buffer[53][7] ) );
  DFFQXL \row1_buffer_reg[52][7]  ( .D(\row1_buffer[53][7] ), .CK(clk), .Q(
        \row1_buffer[52][7] ) );
  DFFQXL \row1_buffer_reg[51][7]  ( .D(\row1_buffer[52][7] ), .CK(clk), .Q(
        \row1_buffer[51][7] ) );
  DFFQXL \row1_buffer_reg[50][7]  ( .D(\row1_buffer[51][7] ), .CK(clk), .Q(
        \row1_buffer[50][7] ) );
  DFFQXL \row1_buffer_reg[49][7]  ( .D(\row1_buffer[50][7] ), .CK(clk), .Q(
        \row1_buffer[49][7] ) );
  DFFQXL \row1_buffer_reg[48][7]  ( .D(\row1_buffer[49][7] ), .CK(clk), .Q(
        \row1_buffer[48][7] ) );
  DFFQXL \row1_buffer_reg[47][7]  ( .D(\row1_buffer[48][7] ), .CK(clk), .Q(
        \row1_buffer[47][7] ) );
  DFFQXL \row1_buffer_reg[46][7]  ( .D(\row1_buffer[47][7] ), .CK(clk), .Q(
        \row1_buffer[46][7] ) );
  DFFQXL \row1_buffer_reg[45][7]  ( .D(\row1_buffer[46][7] ), .CK(clk), .Q(
        \row1_buffer[45][7] ) );
  DFFQXL \row1_buffer_reg[44][7]  ( .D(\row1_buffer[45][7] ), .CK(clk), .Q(
        \row1_buffer[44][7] ) );
  DFFQXL \row1_buffer_reg[43][7]  ( .D(\row1_buffer[44][7] ), .CK(clk), .Q(
        \row1_buffer[43][7] ) );
  DFFQXL \row1_buffer_reg[42][7]  ( .D(\row1_buffer[43][7] ), .CK(clk), .Q(
        \row1_buffer[42][7] ) );
  DFFQXL \row1_buffer_reg[41][7]  ( .D(\row1_buffer[42][7] ), .CK(clk), .Q(
        \row1_buffer[41][7] ) );
  DFFQXL \row1_buffer_reg[40][7]  ( .D(\row1_buffer[41][7] ), .CK(clk), .Q(
        \row1_buffer[40][7] ) );
  DFFQXL \row1_buffer_reg[39][7]  ( .D(\row1_buffer[40][7] ), .CK(clk), .Q(
        \row1_buffer[39][7] ) );
  DFFQXL \row1_buffer_reg[38][7]  ( .D(\row1_buffer[39][7] ), .CK(clk), .Q(
        \row1_buffer[38][7] ) );
  DFFQXL \row1_buffer_reg[37][7]  ( .D(\row1_buffer[38][7] ), .CK(clk), .Q(
        \row1_buffer[37][7] ) );
  DFFQXL \row1_buffer_reg[36][7]  ( .D(\row1_buffer[37][7] ), .CK(clk), .Q(
        \row1_buffer[36][7] ) );
  DFFQXL \row1_buffer_reg[35][7]  ( .D(\row1_buffer[36][7] ), .CK(clk), .Q(
        \row1_buffer[35][7] ) );
  DFFQXL \row1_buffer_reg[34][7]  ( .D(\row1_buffer[35][7] ), .CK(clk), .Q(
        \row1_buffer[34][7] ) );
  DFFQXL \row1_buffer_reg[33][7]  ( .D(\row1_buffer[34][7] ), .CK(clk), .Q(
        \row1_buffer[33][7] ) );
  DFFQXL \row1_buffer_reg[32][7]  ( .D(\row1_buffer[33][7] ), .CK(clk), .Q(
        \row1_buffer[32][7] ) );
  DFFQXL \row1_buffer_reg[31][7]  ( .D(\row1_buffer[32][7] ), .CK(clk), .Q(
        \row1_buffer[31][7] ) );
  DFFQXL \row1_buffer_reg[30][7]  ( .D(\row1_buffer[31][7] ), .CK(clk), .Q(
        \row1_buffer[30][7] ) );
  DFFQXL \row1_buffer_reg[29][7]  ( .D(\row1_buffer[30][7] ), .CK(clk), .Q(
        \row1_buffer[29][7] ) );
  DFFQXL \row1_buffer_reg[28][7]  ( .D(\row1_buffer[29][7] ), .CK(clk), .Q(
        \row1_buffer[28][7] ) );
  DFFQXL \row1_buffer_reg[27][7]  ( .D(\row1_buffer[28][7] ), .CK(clk), .Q(
        \row1_buffer[27][7] ) );
  DFFQXL \row1_buffer_reg[26][7]  ( .D(\row1_buffer[27][7] ), .CK(clk), .Q(
        \row1_buffer[26][7] ) );
  DFFQXL \row1_buffer_reg[25][7]  ( .D(\row1_buffer[26][7] ), .CK(clk), .Q(
        \row1_buffer[25][7] ) );
  DFFQXL \row1_buffer_reg[24][7]  ( .D(\row1_buffer[25][7] ), .CK(clk), .Q(
        \row1_buffer[24][7] ) );
  DFFQXL \row1_buffer_reg[23][7]  ( .D(\row1_buffer[24][7] ), .CK(clk), .Q(
        \row1_buffer[23][7] ) );
  DFFQXL \row1_buffer_reg[22][7]  ( .D(\row1_buffer[23][7] ), .CK(clk), .Q(
        \row1_buffer[22][7] ) );
  DFFQXL \row1_buffer_reg[21][7]  ( .D(\row1_buffer[22][7] ), .CK(clk), .Q(
        \row1_buffer[21][7] ) );
  DFFQXL \row1_buffer_reg[20][7]  ( .D(\row1_buffer[21][7] ), .CK(clk), .Q(
        \row1_buffer[20][7] ) );
  DFFQXL \row1_buffer_reg[19][7]  ( .D(\row1_buffer[20][7] ), .CK(clk), .Q(
        \row1_buffer[19][7] ) );
  DFFQXL \row1_buffer_reg[18][7]  ( .D(\row1_buffer[19][7] ), .CK(clk), .Q(
        \row1_buffer[18][7] ) );
  DFFQXL \row1_buffer_reg[17][7]  ( .D(\row1_buffer[18][7] ), .CK(clk), .Q(
        \row1_buffer[17][7] ) );
  DFFQXL \row1_buffer_reg[16][7]  ( .D(\row1_buffer[17][7] ), .CK(clk), .Q(
        \row1_buffer[16][7] ) );
  DFFQXL \row1_buffer_reg[15][7]  ( .D(\row1_buffer[16][7] ), .CK(clk), .Q(
        \row1_buffer[15][7] ) );
  DFFQXL \row1_buffer_reg[14][7]  ( .D(\row1_buffer[15][7] ), .CK(clk), .Q(
        \row1_buffer[14][7] ) );
  DFFQXL \row1_buffer_reg[13][7]  ( .D(\row1_buffer[14][7] ), .CK(clk), .Q(
        \row1_buffer[13][7] ) );
  DFFQXL \row1_buffer_reg[12][7]  ( .D(\row1_buffer[13][7] ), .CK(clk), .Q(
        \row1_buffer[12][7] ) );
  DFFQXL \row1_buffer_reg[11][7]  ( .D(\row1_buffer[12][7] ), .CK(clk), .Q(
        \row1_buffer[11][7] ) );
  DFFQXL \row1_buffer_reg[10][7]  ( .D(\row1_buffer[11][7] ), .CK(clk), .Q(
        \row1_buffer[10][7] ) );
  DFFQXL \row1_buffer_reg[9][7]  ( .D(\row1_buffer[10][7] ), .CK(clk), .Q(
        \row1_buffer[9][7] ) );
  DFFQXL \row1_buffer_reg[8][7]  ( .D(\row1_buffer[9][7] ), .CK(clk), .Q(
        \row1_buffer[8][7] ) );
  DFFQXL \row1_buffer_reg[7][7]  ( .D(\row1_buffer[8][7] ), .CK(clk), .Q(
        \row1_buffer[7][7] ) );
  DFFQXL \row1_buffer_reg[6][7]  ( .D(\row1_buffer[7][7] ), .CK(clk), .Q(
        \row1_buffer[6][7] ) );
  DFFQXL \row1_buffer_reg[5][7]  ( .D(\row1_buffer[6][7] ), .CK(clk), .Q(
        \row1_buffer[5][7] ) );
  DFFQXL \row1_buffer_reg[4][7]  ( .D(\row1_buffer[5][7] ), .CK(clk), .Q(
        \row1_buffer[4][7] ) );
  DFFQXL \row1_buffer_reg[3][7]  ( .D(\row1_buffer[4][7] ), .CK(clk), .Q(
        \row1_buffer[3][7] ) );
  DFFQXL \row2_buffer_reg[225][6]  ( .D(\row3_buffer[0][6] ), .CK(clk), .Q(
        \row2_buffer[225][6] ) );
  DFFQXL \row2_buffer_reg[224][6]  ( .D(\row2_buffer[225][6] ), .CK(clk), .Q(
        \row2_buffer[224][6] ) );
  DFFQXL \row2_buffer_reg[223][6]  ( .D(\row2_buffer[224][6] ), .CK(clk), .Q(
        \row2_buffer[223][6] ) );
  DFFQXL \row2_buffer_reg[222][6]  ( .D(\row2_buffer[223][6] ), .CK(clk), .Q(
        \row2_buffer[222][6] ) );
  DFFQXL \row2_buffer_reg[221][6]  ( .D(\row2_buffer[222][6] ), .CK(clk), .Q(
        \row2_buffer[221][6] ) );
  DFFQXL \row2_buffer_reg[220][6]  ( .D(\row2_buffer[221][6] ), .CK(clk), .Q(
        \row2_buffer[220][6] ) );
  DFFQXL \row2_buffer_reg[219][6]  ( .D(\row2_buffer[220][6] ), .CK(clk), .Q(
        \row2_buffer[219][6] ) );
  DFFQXL \row2_buffer_reg[218][6]  ( .D(\row2_buffer[219][6] ), .CK(clk), .Q(
        \row2_buffer[218][6] ) );
  DFFQXL \row2_buffer_reg[217][6]  ( .D(\row2_buffer[218][6] ), .CK(clk), .Q(
        \row2_buffer[217][6] ) );
  DFFQXL \row2_buffer_reg[216][6]  ( .D(\row2_buffer[217][6] ), .CK(clk), .Q(
        \row2_buffer[216][6] ) );
  DFFQXL \row2_buffer_reg[215][6]  ( .D(\row2_buffer[216][6] ), .CK(clk), .Q(
        \row2_buffer[215][6] ) );
  DFFQXL \row2_buffer_reg[214][6]  ( .D(\row2_buffer[215][6] ), .CK(clk), .Q(
        \row2_buffer[214][6] ) );
  DFFQXL \row2_buffer_reg[213][6]  ( .D(\row2_buffer[214][6] ), .CK(clk), .Q(
        \row2_buffer[213][6] ) );
  DFFQXL \row2_buffer_reg[212][6]  ( .D(\row2_buffer[213][6] ), .CK(clk), .Q(
        \row2_buffer[212][6] ) );
  DFFQXL \row2_buffer_reg[211][6]  ( .D(\row2_buffer[212][6] ), .CK(clk), .Q(
        \row2_buffer[211][6] ) );
  DFFQXL \row2_buffer_reg[210][6]  ( .D(\row2_buffer[211][6] ), .CK(clk), .Q(
        \row2_buffer[210][6] ) );
  DFFQXL \row2_buffer_reg[209][6]  ( .D(\row2_buffer[210][6] ), .CK(clk), .Q(
        \row2_buffer[209][6] ) );
  DFFQXL \row2_buffer_reg[208][6]  ( .D(\row2_buffer[209][6] ), .CK(clk), .Q(
        \row2_buffer[208][6] ) );
  DFFQXL \row2_buffer_reg[207][6]  ( .D(\row2_buffer[208][6] ), .CK(clk), .Q(
        \row2_buffer[207][6] ) );
  DFFQXL \row2_buffer_reg[206][6]  ( .D(\row2_buffer[207][6] ), .CK(clk), .Q(
        \row2_buffer[206][6] ) );
  DFFQXL \row2_buffer_reg[205][6]  ( .D(\row2_buffer[206][6] ), .CK(clk), .Q(
        \row2_buffer[205][6] ) );
  DFFQXL \row2_buffer_reg[204][6]  ( .D(\row2_buffer[205][6] ), .CK(clk), .Q(
        \row2_buffer[204][6] ) );
  DFFQXL \row2_buffer_reg[203][6]  ( .D(\row2_buffer[204][6] ), .CK(clk), .Q(
        \row2_buffer[203][6] ) );
  DFFQXL \row2_buffer_reg[202][6]  ( .D(\row2_buffer[203][6] ), .CK(clk), .Q(
        \row2_buffer[202][6] ) );
  DFFQXL \row2_buffer_reg[201][6]  ( .D(\row2_buffer[202][6] ), .CK(clk), .Q(
        \row2_buffer[201][6] ) );
  DFFQXL \row2_buffer_reg[200][6]  ( .D(\row2_buffer[201][6] ), .CK(clk), .Q(
        \row2_buffer[200][6] ) );
  DFFQXL \row2_buffer_reg[199][6]  ( .D(\row2_buffer[200][6] ), .CK(clk), .Q(
        \row2_buffer[199][6] ) );
  DFFQXL \row2_buffer_reg[198][6]  ( .D(\row2_buffer[199][6] ), .CK(clk), .Q(
        \row2_buffer[198][6] ) );
  DFFQXL \row2_buffer_reg[197][6]  ( .D(\row2_buffer[198][6] ), .CK(clk), .Q(
        \row2_buffer[197][6] ) );
  DFFQXL \row2_buffer_reg[196][6]  ( .D(\row2_buffer[197][6] ), .CK(clk), .Q(
        \row2_buffer[196][6] ) );
  DFFQXL \row2_buffer_reg[195][6]  ( .D(\row2_buffer[196][6] ), .CK(clk), .Q(
        \row2_buffer[195][6] ) );
  DFFQXL \row2_buffer_reg[194][6]  ( .D(\row2_buffer[195][6] ), .CK(clk), .Q(
        \row2_buffer[194][6] ) );
  DFFQXL \row2_buffer_reg[193][6]  ( .D(\row2_buffer[194][6] ), .CK(clk), .Q(
        \row2_buffer[193][6] ) );
  DFFQXL \row2_buffer_reg[192][6]  ( .D(\row2_buffer[193][6] ), .CK(clk), .Q(
        \row2_buffer[192][6] ) );
  DFFQXL \row2_buffer_reg[191][6]  ( .D(\row2_buffer[192][6] ), .CK(clk), .Q(
        \row2_buffer[191][6] ) );
  DFFQXL \row2_buffer_reg[190][6]  ( .D(\row2_buffer[191][6] ), .CK(clk), .Q(
        \row2_buffer[190][6] ) );
  DFFQXL \row2_buffer_reg[189][6]  ( .D(\row2_buffer[190][6] ), .CK(clk), .Q(
        \row2_buffer[189][6] ) );
  DFFQXL \row2_buffer_reg[188][6]  ( .D(\row2_buffer[189][6] ), .CK(clk), .Q(
        \row2_buffer[188][6] ) );
  DFFQXL \row2_buffer_reg[187][6]  ( .D(\row2_buffer[188][6] ), .CK(clk), .Q(
        \row2_buffer[187][6] ) );
  DFFQXL \row2_buffer_reg[186][6]  ( .D(\row2_buffer[187][6] ), .CK(clk), .Q(
        \row2_buffer[186][6] ) );
  DFFQXL \row2_buffer_reg[185][6]  ( .D(\row2_buffer[186][6] ), .CK(clk), .Q(
        \row2_buffer[185][6] ) );
  DFFQXL \row2_buffer_reg[184][6]  ( .D(\row2_buffer[185][6] ), .CK(clk), .Q(
        \row2_buffer[184][6] ) );
  DFFQXL \row2_buffer_reg[183][6]  ( .D(\row2_buffer[184][6] ), .CK(clk), .Q(
        \row2_buffer[183][6] ) );
  DFFQXL \row2_buffer_reg[182][6]  ( .D(\row2_buffer[183][6] ), .CK(clk), .Q(
        \row2_buffer[182][6] ) );
  DFFQXL \row2_buffer_reg[181][6]  ( .D(\row2_buffer[182][6] ), .CK(clk), .Q(
        \row2_buffer[181][6] ) );
  DFFQXL \row2_buffer_reg[180][6]  ( .D(\row2_buffer[181][6] ), .CK(clk), .Q(
        \row2_buffer[180][6] ) );
  DFFQXL \row2_buffer_reg[179][6]  ( .D(\row2_buffer[180][6] ), .CK(clk), .Q(
        \row2_buffer[179][6] ) );
  DFFQXL \row2_buffer_reg[178][6]  ( .D(\row2_buffer[179][6] ), .CK(clk), .Q(
        \row2_buffer[178][6] ) );
  DFFQXL \row2_buffer_reg[177][6]  ( .D(\row2_buffer[178][6] ), .CK(clk), .Q(
        \row2_buffer[177][6] ) );
  DFFQXL \row2_buffer_reg[176][6]  ( .D(\row2_buffer[177][6] ), .CK(clk), .Q(
        \row2_buffer[176][6] ) );
  DFFQXL \row2_buffer_reg[175][6]  ( .D(\row2_buffer[176][6] ), .CK(clk), .Q(
        \row2_buffer[175][6] ) );
  DFFQXL \row2_buffer_reg[174][6]  ( .D(\row2_buffer[175][6] ), .CK(clk), .Q(
        \row2_buffer[174][6] ) );
  DFFQXL \row2_buffer_reg[173][6]  ( .D(\row2_buffer[174][6] ), .CK(clk), .Q(
        \row2_buffer[173][6] ) );
  DFFQXL \row2_buffer_reg[172][6]  ( .D(\row2_buffer[173][6] ), .CK(clk), .Q(
        \row2_buffer[172][6] ) );
  DFFQXL \row2_buffer_reg[171][6]  ( .D(\row2_buffer[172][6] ), .CK(clk), .Q(
        \row2_buffer[171][6] ) );
  DFFQXL \row2_buffer_reg[170][6]  ( .D(\row2_buffer[171][6] ), .CK(clk), .Q(
        \row2_buffer[170][6] ) );
  DFFQXL \row2_buffer_reg[169][6]  ( .D(\row2_buffer[170][6] ), .CK(clk), .Q(
        \row2_buffer[169][6] ) );
  DFFQXL \row2_buffer_reg[168][6]  ( .D(\row2_buffer[169][6] ), .CK(clk), .Q(
        \row2_buffer[168][6] ) );
  DFFQXL \row2_buffer_reg[167][6]  ( .D(\row2_buffer[168][6] ), .CK(clk), .Q(
        \row2_buffer[167][6] ) );
  DFFQXL \row2_buffer_reg[166][6]  ( .D(\row2_buffer[167][6] ), .CK(clk), .Q(
        \row2_buffer[166][6] ) );
  DFFQXL \row2_buffer_reg[165][6]  ( .D(\row2_buffer[166][6] ), .CK(clk), .Q(
        \row2_buffer[165][6] ) );
  DFFQXL \row2_buffer_reg[164][6]  ( .D(\row2_buffer[165][6] ), .CK(clk), .Q(
        \row2_buffer[164][6] ) );
  DFFQXL \row2_buffer_reg[163][6]  ( .D(\row2_buffer[164][6] ), .CK(clk), .Q(
        \row2_buffer[163][6] ) );
  DFFQXL \row2_buffer_reg[162][6]  ( .D(\row2_buffer[163][6] ), .CK(clk), .Q(
        \row2_buffer[162][6] ) );
  DFFQXL \row2_buffer_reg[161][6]  ( .D(\row2_buffer[162][6] ), .CK(clk), .Q(
        \row2_buffer[161][6] ) );
  DFFQXL \row2_buffer_reg[160][6]  ( .D(\row2_buffer[161][6] ), .CK(clk), .Q(
        \row2_buffer[160][6] ) );
  DFFQXL \row2_buffer_reg[159][6]  ( .D(\row2_buffer[160][6] ), .CK(clk), .Q(
        \row2_buffer[159][6] ) );
  DFFQXL \row2_buffer_reg[158][6]  ( .D(\row2_buffer[159][6] ), .CK(clk), .Q(
        \row2_buffer[158][6] ) );
  DFFQXL \row2_buffer_reg[157][6]  ( .D(\row2_buffer[158][6] ), .CK(clk), .Q(
        \row2_buffer[157][6] ) );
  DFFQXL \row2_buffer_reg[156][6]  ( .D(\row2_buffer[157][6] ), .CK(clk), .Q(
        \row2_buffer[156][6] ) );
  DFFQXL \row2_buffer_reg[155][6]  ( .D(\row2_buffer[156][6] ), .CK(clk), .Q(
        \row2_buffer[155][6] ) );
  DFFQXL \row2_buffer_reg[154][6]  ( .D(\row2_buffer[155][6] ), .CK(clk), .Q(
        \row2_buffer[154][6] ) );
  DFFQXL \row2_buffer_reg[153][6]  ( .D(\row2_buffer[154][6] ), .CK(clk), .Q(
        \row2_buffer[153][6] ) );
  DFFQXL \row2_buffer_reg[152][6]  ( .D(\row2_buffer[153][6] ), .CK(clk), .Q(
        \row2_buffer[152][6] ) );
  DFFQXL \row2_buffer_reg[151][6]  ( .D(\row2_buffer[152][6] ), .CK(clk), .Q(
        \row2_buffer[151][6] ) );
  DFFQXL \row2_buffer_reg[150][6]  ( .D(\row2_buffer[151][6] ), .CK(clk), .Q(
        \row2_buffer[150][6] ) );
  DFFQXL \row2_buffer_reg[149][6]  ( .D(\row2_buffer[150][6] ), .CK(clk), .Q(
        \row2_buffer[149][6] ) );
  DFFQXL \row2_buffer_reg[148][6]  ( .D(\row2_buffer[149][6] ), .CK(clk), .Q(
        \row2_buffer[148][6] ) );
  DFFQXL \row2_buffer_reg[147][6]  ( .D(\row2_buffer[148][6] ), .CK(clk), .Q(
        \row2_buffer[147][6] ) );
  DFFQXL \row2_buffer_reg[146][6]  ( .D(\row2_buffer[147][6] ), .CK(clk), .Q(
        \row2_buffer[146][6] ) );
  DFFQXL \row2_buffer_reg[145][6]  ( .D(\row2_buffer[146][6] ), .CK(clk), .Q(
        \row2_buffer[145][6] ) );
  DFFQXL \row2_buffer_reg[144][6]  ( .D(\row2_buffer[145][6] ), .CK(clk), .Q(
        \row2_buffer[144][6] ) );
  DFFQXL \row2_buffer_reg[143][6]  ( .D(\row2_buffer[144][6] ), .CK(clk), .Q(
        \row2_buffer[143][6] ) );
  DFFQXL \row2_buffer_reg[142][6]  ( .D(\row2_buffer[143][6] ), .CK(clk), .Q(
        \row2_buffer[142][6] ) );
  DFFQXL \row2_buffer_reg[141][6]  ( .D(\row2_buffer[142][6] ), .CK(clk), .Q(
        \row2_buffer[141][6] ) );
  DFFQXL \row2_buffer_reg[140][6]  ( .D(\row2_buffer[141][6] ), .CK(clk), .Q(
        \row2_buffer[140][6] ) );
  DFFQXL \row2_buffer_reg[139][6]  ( .D(\row2_buffer[140][6] ), .CK(clk), .Q(
        \row2_buffer[139][6] ) );
  DFFQXL \row2_buffer_reg[138][6]  ( .D(\row2_buffer[139][6] ), .CK(clk), .Q(
        \row2_buffer[138][6] ) );
  DFFQXL \row2_buffer_reg[137][6]  ( .D(\row2_buffer[138][6] ), .CK(clk), .Q(
        \row2_buffer[137][6] ) );
  DFFQXL \row2_buffer_reg[136][6]  ( .D(\row2_buffer[137][6] ), .CK(clk), .Q(
        \row2_buffer[136][6] ) );
  DFFQXL \row2_buffer_reg[135][6]  ( .D(\row2_buffer[136][6] ), .CK(clk), .Q(
        \row2_buffer[135][6] ) );
  DFFQXL \row2_buffer_reg[134][6]  ( .D(\row2_buffer[135][6] ), .CK(clk), .Q(
        \row2_buffer[134][6] ) );
  DFFQXL \row2_buffer_reg[133][6]  ( .D(\row2_buffer[134][6] ), .CK(clk), .Q(
        \row2_buffer[133][6] ) );
  DFFQXL \row2_buffer_reg[132][6]  ( .D(\row2_buffer[133][6] ), .CK(clk), .Q(
        \row2_buffer[132][6] ) );
  DFFQXL \row2_buffer_reg[131][6]  ( .D(\row2_buffer[132][6] ), .CK(clk), .Q(
        \row2_buffer[131][6] ) );
  DFFQXL \row2_buffer_reg[130][6]  ( .D(\row2_buffer[131][6] ), .CK(clk), .Q(
        \row2_buffer[130][6] ) );
  DFFQXL \row2_buffer_reg[129][6]  ( .D(\row2_buffer[130][6] ), .CK(clk), .Q(
        \row2_buffer[129][6] ) );
  DFFQXL \row2_buffer_reg[128][6]  ( .D(\row2_buffer[129][6] ), .CK(clk), .Q(
        \row2_buffer[128][6] ) );
  DFFQXL \row2_buffer_reg[127][6]  ( .D(\row2_buffer[128][6] ), .CK(clk), .Q(
        \row2_buffer[127][6] ) );
  DFFQXL \row2_buffer_reg[126][6]  ( .D(\row2_buffer[127][6] ), .CK(clk), .Q(
        \row2_buffer[126][6] ) );
  DFFQXL \row2_buffer_reg[125][6]  ( .D(\row2_buffer[126][6] ), .CK(clk), .Q(
        \row2_buffer[125][6] ) );
  DFFQXL \row2_buffer_reg[124][6]  ( .D(\row2_buffer[125][6] ), .CK(clk), .Q(
        \row2_buffer[124][6] ) );
  DFFQXL \row2_buffer_reg[123][6]  ( .D(\row2_buffer[124][6] ), .CK(clk), .Q(
        \row2_buffer[123][6] ) );
  DFFQXL \row2_buffer_reg[122][6]  ( .D(\row2_buffer[123][6] ), .CK(clk), .Q(
        \row2_buffer[122][6] ) );
  DFFQXL \row2_buffer_reg[121][6]  ( .D(\row2_buffer[122][6] ), .CK(clk), .Q(
        \row2_buffer[121][6] ) );
  DFFQXL \row2_buffer_reg[120][6]  ( .D(\row2_buffer[121][6] ), .CK(clk), .Q(
        \row2_buffer[120][6] ) );
  DFFQXL \row2_buffer_reg[119][6]  ( .D(\row2_buffer[120][6] ), .CK(clk), .Q(
        \row2_buffer[119][6] ) );
  DFFQXL \row2_buffer_reg[118][6]  ( .D(\row2_buffer[119][6] ), .CK(clk), .Q(
        \row2_buffer[118][6] ) );
  DFFQXL \row2_buffer_reg[117][6]  ( .D(\row2_buffer[118][6] ), .CK(clk), .Q(
        \row2_buffer[117][6] ) );
  DFFQXL \row2_buffer_reg[116][6]  ( .D(\row2_buffer[117][6] ), .CK(clk), .Q(
        \row2_buffer[116][6] ) );
  DFFQXL \row2_buffer_reg[115][6]  ( .D(\row2_buffer[116][6] ), .CK(clk), .Q(
        \row2_buffer[115][6] ) );
  DFFQXL \row2_buffer_reg[114][6]  ( .D(\row2_buffer[115][6] ), .CK(clk), .Q(
        \row2_buffer[114][6] ) );
  DFFQXL \row2_buffer_reg[113][6]  ( .D(\row2_buffer[114][6] ), .CK(clk), .Q(
        \row2_buffer[113][6] ) );
  DFFQXL \row2_buffer_reg[112][6]  ( .D(\row2_buffer[113][6] ), .CK(clk), .Q(
        \row2_buffer[112][6] ) );
  DFFQXL \row2_buffer_reg[111][6]  ( .D(\row2_buffer[112][6] ), .CK(clk), .Q(
        \row2_buffer[111][6] ) );
  DFFQXL \row2_buffer_reg[110][6]  ( .D(\row2_buffer[111][6] ), .CK(clk), .Q(
        \row2_buffer[110][6] ) );
  DFFQXL \row2_buffer_reg[109][6]  ( .D(\row2_buffer[110][6] ), .CK(clk), .Q(
        \row2_buffer[109][6] ) );
  DFFQXL \row2_buffer_reg[108][6]  ( .D(\row2_buffer[109][6] ), .CK(clk), .Q(
        \row2_buffer[108][6] ) );
  DFFQXL \row2_buffer_reg[107][6]  ( .D(\row2_buffer[108][6] ), .CK(clk), .Q(
        \row2_buffer[107][6] ) );
  DFFQXL \row2_buffer_reg[106][6]  ( .D(\row2_buffer[107][6] ), .CK(clk), .Q(
        \row2_buffer[106][6] ) );
  DFFQXL \row2_buffer_reg[105][6]  ( .D(\row2_buffer[106][6] ), .CK(clk), .Q(
        \row2_buffer[105][6] ) );
  DFFQXL \row2_buffer_reg[104][6]  ( .D(\row2_buffer[105][6] ), .CK(clk), .Q(
        \row2_buffer[104][6] ) );
  DFFQXL \row2_buffer_reg[103][6]  ( .D(\row2_buffer[104][6] ), .CK(clk), .Q(
        \row2_buffer[103][6] ) );
  DFFQXL \row2_buffer_reg[102][6]  ( .D(\row2_buffer[103][6] ), .CK(clk), .Q(
        \row2_buffer[102][6] ) );
  DFFQXL \row2_buffer_reg[101][6]  ( .D(\row2_buffer[102][6] ), .CK(clk), .Q(
        \row2_buffer[101][6] ) );
  DFFQXL \row2_buffer_reg[100][6]  ( .D(\row2_buffer[101][6] ), .CK(clk), .Q(
        \row2_buffer[100][6] ) );
  DFFQXL \row2_buffer_reg[99][6]  ( .D(\row2_buffer[100][6] ), .CK(clk), .Q(
        \row2_buffer[99][6] ) );
  DFFQXL \row2_buffer_reg[98][6]  ( .D(\row2_buffer[99][6] ), .CK(clk), .Q(
        \row2_buffer[98][6] ) );
  DFFQXL \row2_buffer_reg[97][6]  ( .D(\row2_buffer[98][6] ), .CK(clk), .Q(
        \row2_buffer[97][6] ) );
  DFFQXL \row2_buffer_reg[96][6]  ( .D(\row2_buffer[97][6] ), .CK(clk), .Q(
        \row2_buffer[96][6] ) );
  DFFQXL \row2_buffer_reg[95][6]  ( .D(\row2_buffer[96][6] ), .CK(clk), .Q(
        \row2_buffer[95][6] ) );
  DFFQXL \row2_buffer_reg[94][6]  ( .D(\row2_buffer[95][6] ), .CK(clk), .Q(
        \row2_buffer[94][6] ) );
  DFFQXL \row2_buffer_reg[93][6]  ( .D(\row2_buffer[94][6] ), .CK(clk), .Q(
        \row2_buffer[93][6] ) );
  DFFQXL \row2_buffer_reg[92][6]  ( .D(\row2_buffer[93][6] ), .CK(clk), .Q(
        \row2_buffer[92][6] ) );
  DFFQXL \row2_buffer_reg[91][6]  ( .D(\row2_buffer[92][6] ), .CK(clk), .Q(
        \row2_buffer[91][6] ) );
  DFFQXL \row2_buffer_reg[90][6]  ( .D(\row2_buffer[91][6] ), .CK(clk), .Q(
        \row2_buffer[90][6] ) );
  DFFQXL \row2_buffer_reg[89][6]  ( .D(\row2_buffer[90][6] ), .CK(clk), .Q(
        \row2_buffer[89][6] ) );
  DFFQXL \row2_buffer_reg[88][6]  ( .D(\row2_buffer[89][6] ), .CK(clk), .Q(
        \row2_buffer[88][6] ) );
  DFFQXL \row2_buffer_reg[87][6]  ( .D(\row2_buffer[88][6] ), .CK(clk), .Q(
        \row2_buffer[87][6] ) );
  DFFQXL \row2_buffer_reg[86][6]  ( .D(\row2_buffer[87][6] ), .CK(clk), .Q(
        \row2_buffer[86][6] ) );
  DFFQXL \row2_buffer_reg[85][6]  ( .D(\row2_buffer[86][6] ), .CK(clk), .Q(
        \row2_buffer[85][6] ) );
  DFFQXL \row2_buffer_reg[84][6]  ( .D(\row2_buffer[85][6] ), .CK(clk), .Q(
        \row2_buffer[84][6] ) );
  DFFQXL \row2_buffer_reg[83][6]  ( .D(\row2_buffer[84][6] ), .CK(clk), .Q(
        \row2_buffer[83][6] ) );
  DFFQXL \row2_buffer_reg[82][6]  ( .D(\row2_buffer[83][6] ), .CK(clk), .Q(
        \row2_buffer[82][6] ) );
  DFFQXL \row2_buffer_reg[81][6]  ( .D(\row2_buffer[82][6] ), .CK(clk), .Q(
        \row2_buffer[81][6] ) );
  DFFQXL \row2_buffer_reg[80][6]  ( .D(\row2_buffer[81][6] ), .CK(clk), .Q(
        \row2_buffer[80][6] ) );
  DFFQXL \row2_buffer_reg[79][6]  ( .D(\row2_buffer[80][6] ), .CK(clk), .Q(
        \row2_buffer[79][6] ) );
  DFFQXL \row2_buffer_reg[78][6]  ( .D(\row2_buffer[79][6] ), .CK(clk), .Q(
        \row2_buffer[78][6] ) );
  DFFQXL \row2_buffer_reg[77][6]  ( .D(\row2_buffer[78][6] ), .CK(clk), .Q(
        \row2_buffer[77][6] ) );
  DFFQXL \row2_buffer_reg[76][6]  ( .D(\row2_buffer[77][6] ), .CK(clk), .Q(
        \row2_buffer[76][6] ) );
  DFFQXL \row2_buffer_reg[75][6]  ( .D(\row2_buffer[76][6] ), .CK(clk), .Q(
        \row2_buffer[75][6] ) );
  DFFQXL \row2_buffer_reg[74][6]  ( .D(\row2_buffer[75][6] ), .CK(clk), .Q(
        \row2_buffer[74][6] ) );
  DFFQXL \row2_buffer_reg[73][6]  ( .D(\row2_buffer[74][6] ), .CK(clk), .Q(
        \row2_buffer[73][6] ) );
  DFFQXL \row2_buffer_reg[72][6]  ( .D(\row2_buffer[73][6] ), .CK(clk), .Q(
        \row2_buffer[72][6] ) );
  DFFQXL \row2_buffer_reg[71][6]  ( .D(\row2_buffer[72][6] ), .CK(clk), .Q(
        \row2_buffer[71][6] ) );
  DFFQXL \row2_buffer_reg[70][6]  ( .D(\row2_buffer[71][6] ), .CK(clk), .Q(
        \row2_buffer[70][6] ) );
  DFFQXL \row2_buffer_reg[69][6]  ( .D(\row2_buffer[70][6] ), .CK(clk), .Q(
        \row2_buffer[69][6] ) );
  DFFQXL \row2_buffer_reg[68][6]  ( .D(\row2_buffer[69][6] ), .CK(clk), .Q(
        \row2_buffer[68][6] ) );
  DFFQXL \row2_buffer_reg[67][6]  ( .D(\row2_buffer[68][6] ), .CK(clk), .Q(
        \row2_buffer[67][6] ) );
  DFFQXL \row2_buffer_reg[66][6]  ( .D(\row2_buffer[67][6] ), .CK(clk), .Q(
        \row2_buffer[66][6] ) );
  DFFQXL \row2_buffer_reg[65][6]  ( .D(\row2_buffer[66][6] ), .CK(clk), .Q(
        \row2_buffer[65][6] ) );
  DFFQXL \row2_buffer_reg[64][6]  ( .D(\row2_buffer[65][6] ), .CK(clk), .Q(
        \row2_buffer[64][6] ) );
  DFFQXL \row2_buffer_reg[63][6]  ( .D(\row2_buffer[64][6] ), .CK(clk), .Q(
        \row2_buffer[63][6] ) );
  DFFQXL \row2_buffer_reg[62][6]  ( .D(\row2_buffer[63][6] ), .CK(clk), .Q(
        \row2_buffer[62][6] ) );
  DFFQXL \row2_buffer_reg[61][6]  ( .D(\row2_buffer[62][6] ), .CK(clk), .Q(
        \row2_buffer[61][6] ) );
  DFFQXL \row2_buffer_reg[60][6]  ( .D(\row2_buffer[61][6] ), .CK(clk), .Q(
        \row2_buffer[60][6] ) );
  DFFQXL \row2_buffer_reg[59][6]  ( .D(\row2_buffer[60][6] ), .CK(clk), .Q(
        \row2_buffer[59][6] ) );
  DFFQXL \row2_buffer_reg[58][6]  ( .D(\row2_buffer[59][6] ), .CK(clk), .Q(
        \row2_buffer[58][6] ) );
  DFFQXL \row2_buffer_reg[57][6]  ( .D(\row2_buffer[58][6] ), .CK(clk), .Q(
        \row2_buffer[57][6] ) );
  DFFQXL \row2_buffer_reg[56][6]  ( .D(\row2_buffer[57][6] ), .CK(clk), .Q(
        \row2_buffer[56][6] ) );
  DFFQXL \row2_buffer_reg[55][6]  ( .D(\row2_buffer[56][6] ), .CK(clk), .Q(
        \row2_buffer[55][6] ) );
  DFFQXL \row2_buffer_reg[54][6]  ( .D(\row2_buffer[55][6] ), .CK(clk), .Q(
        \row2_buffer[54][6] ) );
  DFFQXL \row2_buffer_reg[53][6]  ( .D(\row2_buffer[54][6] ), .CK(clk), .Q(
        \row2_buffer[53][6] ) );
  DFFQXL \row2_buffer_reg[52][6]  ( .D(\row2_buffer[53][6] ), .CK(clk), .Q(
        \row2_buffer[52][6] ) );
  DFFQXL \row2_buffer_reg[51][6]  ( .D(\row2_buffer[52][6] ), .CK(clk), .Q(
        \row2_buffer[51][6] ) );
  DFFQXL \row2_buffer_reg[50][6]  ( .D(\row2_buffer[51][6] ), .CK(clk), .Q(
        \row2_buffer[50][6] ) );
  DFFQXL \row2_buffer_reg[49][6]  ( .D(\row2_buffer[50][6] ), .CK(clk), .Q(
        \row2_buffer[49][6] ) );
  DFFQXL \row2_buffer_reg[48][6]  ( .D(\row2_buffer[49][6] ), .CK(clk), .Q(
        \row2_buffer[48][6] ) );
  DFFQXL \row2_buffer_reg[47][6]  ( .D(\row2_buffer[48][6] ), .CK(clk), .Q(
        \row2_buffer[47][6] ) );
  DFFQXL \row2_buffer_reg[46][6]  ( .D(\row2_buffer[47][6] ), .CK(clk), .Q(
        \row2_buffer[46][6] ) );
  DFFQXL \row2_buffer_reg[45][6]  ( .D(\row2_buffer[46][6] ), .CK(clk), .Q(
        \row2_buffer[45][6] ) );
  DFFQXL \row2_buffer_reg[44][6]  ( .D(\row2_buffer[45][6] ), .CK(clk), .Q(
        \row2_buffer[44][6] ) );
  DFFQXL \row2_buffer_reg[43][6]  ( .D(\row2_buffer[44][6] ), .CK(clk), .Q(
        \row2_buffer[43][6] ) );
  DFFQXL \row2_buffer_reg[42][6]  ( .D(\row2_buffer[43][6] ), .CK(clk), .Q(
        \row2_buffer[42][6] ) );
  DFFQXL \row2_buffer_reg[41][6]  ( .D(\row2_buffer[42][6] ), .CK(clk), .Q(
        \row2_buffer[41][6] ) );
  DFFQXL \row2_buffer_reg[40][6]  ( .D(\row2_buffer[41][6] ), .CK(clk), .Q(
        \row2_buffer[40][6] ) );
  DFFQXL \row2_buffer_reg[39][6]  ( .D(\row2_buffer[40][6] ), .CK(clk), .Q(
        \row2_buffer[39][6] ) );
  DFFQXL \row2_buffer_reg[38][6]  ( .D(\row2_buffer[39][6] ), .CK(clk), .Q(
        \row2_buffer[38][6] ) );
  DFFQXL \row2_buffer_reg[37][6]  ( .D(\row2_buffer[38][6] ), .CK(clk), .Q(
        \row2_buffer[37][6] ) );
  DFFQXL \row2_buffer_reg[36][6]  ( .D(\row2_buffer[37][6] ), .CK(clk), .Q(
        \row2_buffer[36][6] ) );
  DFFQXL \row2_buffer_reg[35][6]  ( .D(\row2_buffer[36][6] ), .CK(clk), .Q(
        \row2_buffer[35][6] ) );
  DFFQXL \row2_buffer_reg[34][6]  ( .D(\row2_buffer[35][6] ), .CK(clk), .Q(
        \row2_buffer[34][6] ) );
  DFFQXL \row2_buffer_reg[33][6]  ( .D(\row2_buffer[34][6] ), .CK(clk), .Q(
        \row2_buffer[33][6] ) );
  DFFQXL \row2_buffer_reg[32][6]  ( .D(\row2_buffer[33][6] ), .CK(clk), .Q(
        \row2_buffer[32][6] ) );
  DFFQXL \row2_buffer_reg[31][6]  ( .D(\row2_buffer[32][6] ), .CK(clk), .Q(
        \row2_buffer[31][6] ) );
  DFFQXL \row2_buffer_reg[30][6]  ( .D(\row2_buffer[31][6] ), .CK(clk), .Q(
        \row2_buffer[30][6] ) );
  DFFQXL \row2_buffer_reg[29][6]  ( .D(\row2_buffer[30][6] ), .CK(clk), .Q(
        \row2_buffer[29][6] ) );
  DFFQXL \row2_buffer_reg[28][6]  ( .D(\row2_buffer[29][6] ), .CK(clk), .Q(
        \row2_buffer[28][6] ) );
  DFFQXL \row2_buffer_reg[27][6]  ( .D(\row2_buffer[28][6] ), .CK(clk), .Q(
        \row2_buffer[27][6] ) );
  DFFQXL \row2_buffer_reg[26][6]  ( .D(\row2_buffer[27][6] ), .CK(clk), .Q(
        \row2_buffer[26][6] ) );
  DFFQXL \row2_buffer_reg[25][6]  ( .D(\row2_buffer[26][6] ), .CK(clk), .Q(
        \row2_buffer[25][6] ) );
  DFFQXL \row2_buffer_reg[24][6]  ( .D(\row2_buffer[25][6] ), .CK(clk), .Q(
        \row2_buffer[24][6] ) );
  DFFQXL \row2_buffer_reg[23][6]  ( .D(\row2_buffer[24][6] ), .CK(clk), .Q(
        \row2_buffer[23][6] ) );
  DFFQXL \row2_buffer_reg[22][6]  ( .D(\row2_buffer[23][6] ), .CK(clk), .Q(
        \row2_buffer[22][6] ) );
  DFFQXL \row2_buffer_reg[21][6]  ( .D(\row2_buffer[22][6] ), .CK(clk), .Q(
        \row2_buffer[21][6] ) );
  DFFQXL \row2_buffer_reg[20][6]  ( .D(\row2_buffer[21][6] ), .CK(clk), .Q(
        \row2_buffer[20][6] ) );
  DFFQXL \row2_buffer_reg[19][6]  ( .D(\row2_buffer[20][6] ), .CK(clk), .Q(
        \row2_buffer[19][6] ) );
  DFFQXL \row2_buffer_reg[18][6]  ( .D(\row2_buffer[19][6] ), .CK(clk), .Q(
        \row2_buffer[18][6] ) );
  DFFQXL \row2_buffer_reg[17][6]  ( .D(\row2_buffer[18][6] ), .CK(clk), .Q(
        \row2_buffer[17][6] ) );
  DFFQXL \row2_buffer_reg[16][6]  ( .D(\row2_buffer[17][6] ), .CK(clk), .Q(
        \row2_buffer[16][6] ) );
  DFFQXL \row2_buffer_reg[15][6]  ( .D(\row2_buffer[16][6] ), .CK(clk), .Q(
        \row2_buffer[15][6] ) );
  DFFQXL \row2_buffer_reg[14][6]  ( .D(\row2_buffer[15][6] ), .CK(clk), .Q(
        \row2_buffer[14][6] ) );
  DFFQXL \row2_buffer_reg[13][6]  ( .D(\row2_buffer[14][6] ), .CK(clk), .Q(
        \row2_buffer[13][6] ) );
  DFFQXL \row2_buffer_reg[12][6]  ( .D(\row2_buffer[13][6] ), .CK(clk), .Q(
        \row2_buffer[12][6] ) );
  DFFQXL \row2_buffer_reg[11][6]  ( .D(\row2_buffer[12][6] ), .CK(clk), .Q(
        \row2_buffer[11][6] ) );
  DFFQXL \row2_buffer_reg[10][6]  ( .D(\row2_buffer[11][6] ), .CK(clk), .Q(
        \row2_buffer[10][6] ) );
  DFFQXL \row2_buffer_reg[9][6]  ( .D(\row2_buffer[10][6] ), .CK(clk), .Q(
        \row2_buffer[9][6] ) );
  DFFQXL \row2_buffer_reg[8][6]  ( .D(\row2_buffer[9][6] ), .CK(clk), .Q(
        \row2_buffer[8][6] ) );
  DFFQXL \row2_buffer_reg[7][6]  ( .D(\row2_buffer[8][6] ), .CK(clk), .Q(
        \row2_buffer[7][6] ) );
  DFFQXL \row2_buffer_reg[6][6]  ( .D(\row2_buffer[7][6] ), .CK(clk), .Q(
        \row2_buffer[6][6] ) );
  DFFQXL \row2_buffer_reg[5][6]  ( .D(\row2_buffer[6][6] ), .CK(clk), .Q(
        \row2_buffer[5][6] ) );
  DFFQXL \row2_buffer_reg[4][6]  ( .D(\row2_buffer[5][6] ), .CK(clk), .Q(
        \row2_buffer[4][6] ) );
  DFFQXL \row2_buffer_reg[3][6]  ( .D(\row2_buffer[4][6] ), .CK(clk), .Q(
        \row2_buffer[3][6] ) );
  DFFQXL \row1_buffer_reg[225][6]  ( .D(\row2_buffer[0][6] ), .CK(clk), .Q(
        \row1_buffer[225][6] ) );
  DFFQXL \row1_buffer_reg[224][6]  ( .D(\row1_buffer[225][6] ), .CK(clk), .Q(
        \row1_buffer[224][6] ) );
  DFFQXL \row1_buffer_reg[223][6]  ( .D(\row1_buffer[224][6] ), .CK(clk), .Q(
        \row1_buffer[223][6] ) );
  DFFQXL \row1_buffer_reg[222][6]  ( .D(\row1_buffer[223][6] ), .CK(clk), .Q(
        \row1_buffer[222][6] ) );
  DFFQXL \row1_buffer_reg[221][6]  ( .D(\row1_buffer[222][6] ), .CK(clk), .Q(
        \row1_buffer[221][6] ) );
  DFFQXL \row1_buffer_reg[220][6]  ( .D(\row1_buffer[221][6] ), .CK(clk), .Q(
        \row1_buffer[220][6] ) );
  DFFQXL \row1_buffer_reg[219][6]  ( .D(\row1_buffer[220][6] ), .CK(clk), .Q(
        \row1_buffer[219][6] ) );
  DFFQXL \row1_buffer_reg[218][6]  ( .D(\row1_buffer[219][6] ), .CK(clk), .Q(
        \row1_buffer[218][6] ) );
  DFFQXL \row1_buffer_reg[217][6]  ( .D(\row1_buffer[218][6] ), .CK(clk), .Q(
        \row1_buffer[217][6] ) );
  DFFQXL \row1_buffer_reg[216][6]  ( .D(\row1_buffer[217][6] ), .CK(clk), .Q(
        \row1_buffer[216][6] ) );
  DFFQXL \row1_buffer_reg[215][6]  ( .D(\row1_buffer[216][6] ), .CK(clk), .Q(
        \row1_buffer[215][6] ) );
  DFFQXL \row1_buffer_reg[214][6]  ( .D(\row1_buffer[215][6] ), .CK(clk), .Q(
        \row1_buffer[214][6] ) );
  DFFQXL \row1_buffer_reg[213][6]  ( .D(\row1_buffer[214][6] ), .CK(clk), .Q(
        \row1_buffer[213][6] ) );
  DFFQXL \row1_buffer_reg[212][6]  ( .D(\row1_buffer[213][6] ), .CK(clk), .Q(
        \row1_buffer[212][6] ) );
  DFFQXL \row1_buffer_reg[211][6]  ( .D(\row1_buffer[212][6] ), .CK(clk), .Q(
        \row1_buffer[211][6] ) );
  DFFQXL \row1_buffer_reg[210][6]  ( .D(\row1_buffer[211][6] ), .CK(clk), .Q(
        \row1_buffer[210][6] ) );
  DFFQXL \row1_buffer_reg[209][6]  ( .D(\row1_buffer[210][6] ), .CK(clk), .Q(
        \row1_buffer[209][6] ) );
  DFFQXL \row1_buffer_reg[208][6]  ( .D(\row1_buffer[209][6] ), .CK(clk), .Q(
        \row1_buffer[208][6] ) );
  DFFQXL \row1_buffer_reg[207][6]  ( .D(\row1_buffer[208][6] ), .CK(clk), .Q(
        \row1_buffer[207][6] ) );
  DFFQXL \row1_buffer_reg[206][6]  ( .D(\row1_buffer[207][6] ), .CK(clk), .Q(
        \row1_buffer[206][6] ) );
  DFFQXL \row1_buffer_reg[205][6]  ( .D(\row1_buffer[206][6] ), .CK(clk), .Q(
        \row1_buffer[205][6] ) );
  DFFQXL \row1_buffer_reg[204][6]  ( .D(\row1_buffer[205][6] ), .CK(clk), .Q(
        \row1_buffer[204][6] ) );
  DFFQXL \row1_buffer_reg[203][6]  ( .D(\row1_buffer[204][6] ), .CK(clk), .Q(
        \row1_buffer[203][6] ) );
  DFFQXL \row1_buffer_reg[202][6]  ( .D(\row1_buffer[203][6] ), .CK(clk), .Q(
        \row1_buffer[202][6] ) );
  DFFQXL \row1_buffer_reg[201][6]  ( .D(\row1_buffer[202][6] ), .CK(clk), .Q(
        \row1_buffer[201][6] ) );
  DFFQXL \row1_buffer_reg[200][6]  ( .D(\row1_buffer[201][6] ), .CK(clk), .Q(
        \row1_buffer[200][6] ) );
  DFFQXL \row1_buffer_reg[199][6]  ( .D(\row1_buffer[200][6] ), .CK(clk), .Q(
        \row1_buffer[199][6] ) );
  DFFQXL \row1_buffer_reg[198][6]  ( .D(\row1_buffer[199][6] ), .CK(clk), .Q(
        \row1_buffer[198][6] ) );
  DFFQXL \row1_buffer_reg[197][6]  ( .D(\row1_buffer[198][6] ), .CK(clk), .Q(
        \row1_buffer[197][6] ) );
  DFFQXL \row1_buffer_reg[196][6]  ( .D(\row1_buffer[197][6] ), .CK(clk), .Q(
        \row1_buffer[196][6] ) );
  DFFQXL \row1_buffer_reg[195][6]  ( .D(\row1_buffer[196][6] ), .CK(clk), .Q(
        \row1_buffer[195][6] ) );
  DFFQXL \row1_buffer_reg[194][6]  ( .D(\row1_buffer[195][6] ), .CK(clk), .Q(
        \row1_buffer[194][6] ) );
  DFFQXL \row1_buffer_reg[193][6]  ( .D(\row1_buffer[194][6] ), .CK(clk), .Q(
        \row1_buffer[193][6] ) );
  DFFQXL \row1_buffer_reg[192][6]  ( .D(\row1_buffer[193][6] ), .CK(clk), .Q(
        \row1_buffer[192][6] ) );
  DFFQXL \row1_buffer_reg[191][6]  ( .D(\row1_buffer[192][6] ), .CK(clk), .Q(
        \row1_buffer[191][6] ) );
  DFFQXL \row1_buffer_reg[190][6]  ( .D(\row1_buffer[191][6] ), .CK(clk), .Q(
        \row1_buffer[190][6] ) );
  DFFQXL \row1_buffer_reg[189][6]  ( .D(\row1_buffer[190][6] ), .CK(clk), .Q(
        \row1_buffer[189][6] ) );
  DFFQXL \row1_buffer_reg[188][6]  ( .D(\row1_buffer[189][6] ), .CK(clk), .Q(
        \row1_buffer[188][6] ) );
  DFFQXL \row1_buffer_reg[187][6]  ( .D(\row1_buffer[188][6] ), .CK(clk), .Q(
        \row1_buffer[187][6] ) );
  DFFQXL \row1_buffer_reg[186][6]  ( .D(\row1_buffer[187][6] ), .CK(clk), .Q(
        \row1_buffer[186][6] ) );
  DFFQXL \row1_buffer_reg[185][6]  ( .D(\row1_buffer[186][6] ), .CK(clk), .Q(
        \row1_buffer[185][6] ) );
  DFFQXL \row1_buffer_reg[184][6]  ( .D(\row1_buffer[185][6] ), .CK(clk), .Q(
        \row1_buffer[184][6] ) );
  DFFQXL \row1_buffer_reg[183][6]  ( .D(\row1_buffer[184][6] ), .CK(clk), .Q(
        \row1_buffer[183][6] ) );
  DFFQXL \row1_buffer_reg[182][6]  ( .D(\row1_buffer[183][6] ), .CK(clk), .Q(
        \row1_buffer[182][6] ) );
  DFFQXL \row1_buffer_reg[181][6]  ( .D(\row1_buffer[182][6] ), .CK(clk), .Q(
        \row1_buffer[181][6] ) );
  DFFQXL \row1_buffer_reg[180][6]  ( .D(\row1_buffer[181][6] ), .CK(clk), .Q(
        \row1_buffer[180][6] ) );
  DFFQXL \row1_buffer_reg[179][6]  ( .D(\row1_buffer[180][6] ), .CK(clk), .Q(
        \row1_buffer[179][6] ) );
  DFFQXL \row1_buffer_reg[178][6]  ( .D(\row1_buffer[179][6] ), .CK(clk), .Q(
        \row1_buffer[178][6] ) );
  DFFQXL \row1_buffer_reg[177][6]  ( .D(\row1_buffer[178][6] ), .CK(clk), .Q(
        \row1_buffer[177][6] ) );
  DFFQXL \row1_buffer_reg[176][6]  ( .D(\row1_buffer[177][6] ), .CK(clk), .Q(
        \row1_buffer[176][6] ) );
  DFFQXL \row1_buffer_reg[175][6]  ( .D(\row1_buffer[176][6] ), .CK(clk), .Q(
        \row1_buffer[175][6] ) );
  DFFQXL \row1_buffer_reg[174][6]  ( .D(\row1_buffer[175][6] ), .CK(clk), .Q(
        \row1_buffer[174][6] ) );
  DFFQXL \row1_buffer_reg[173][6]  ( .D(\row1_buffer[174][6] ), .CK(clk), .Q(
        \row1_buffer[173][6] ) );
  DFFQXL \row1_buffer_reg[172][6]  ( .D(\row1_buffer[173][6] ), .CK(clk), .Q(
        \row1_buffer[172][6] ) );
  DFFQXL \row1_buffer_reg[171][6]  ( .D(\row1_buffer[172][6] ), .CK(clk), .Q(
        \row1_buffer[171][6] ) );
  DFFQXL \row1_buffer_reg[170][6]  ( .D(\row1_buffer[171][6] ), .CK(clk), .Q(
        \row1_buffer[170][6] ) );
  DFFQXL \row1_buffer_reg[169][6]  ( .D(\row1_buffer[170][6] ), .CK(clk), .Q(
        \row1_buffer[169][6] ) );
  DFFQXL \row1_buffer_reg[168][6]  ( .D(\row1_buffer[169][6] ), .CK(clk), .Q(
        \row1_buffer[168][6] ) );
  DFFQXL \row1_buffer_reg[167][6]  ( .D(\row1_buffer[168][6] ), .CK(clk), .Q(
        \row1_buffer[167][6] ) );
  DFFQXL \row1_buffer_reg[166][6]  ( .D(\row1_buffer[167][6] ), .CK(clk), .Q(
        \row1_buffer[166][6] ) );
  DFFQXL \row1_buffer_reg[165][6]  ( .D(\row1_buffer[166][6] ), .CK(clk), .Q(
        \row1_buffer[165][6] ) );
  DFFQXL \row1_buffer_reg[164][6]  ( .D(\row1_buffer[165][6] ), .CK(clk), .Q(
        \row1_buffer[164][6] ) );
  DFFQXL \row1_buffer_reg[163][6]  ( .D(\row1_buffer[164][6] ), .CK(clk), .Q(
        \row1_buffer[163][6] ) );
  DFFQXL \row1_buffer_reg[162][6]  ( .D(\row1_buffer[163][6] ), .CK(clk), .Q(
        \row1_buffer[162][6] ) );
  DFFQXL \row1_buffer_reg[161][6]  ( .D(\row1_buffer[162][6] ), .CK(clk), .Q(
        \row1_buffer[161][6] ) );
  DFFQXL \row1_buffer_reg[160][6]  ( .D(\row1_buffer[161][6] ), .CK(clk), .Q(
        \row1_buffer[160][6] ) );
  DFFQXL \row1_buffer_reg[159][6]  ( .D(\row1_buffer[160][6] ), .CK(clk), .Q(
        \row1_buffer[159][6] ) );
  DFFQXL \row1_buffer_reg[158][6]  ( .D(\row1_buffer[159][6] ), .CK(clk), .Q(
        \row1_buffer[158][6] ) );
  DFFQXL \row1_buffer_reg[157][6]  ( .D(\row1_buffer[158][6] ), .CK(clk), .Q(
        \row1_buffer[157][6] ) );
  DFFQXL \row1_buffer_reg[156][6]  ( .D(\row1_buffer[157][6] ), .CK(clk), .Q(
        \row1_buffer[156][6] ) );
  DFFQXL \row1_buffer_reg[155][6]  ( .D(\row1_buffer[156][6] ), .CK(clk), .Q(
        \row1_buffer[155][6] ) );
  DFFQXL \row1_buffer_reg[154][6]  ( .D(\row1_buffer[155][6] ), .CK(clk), .Q(
        \row1_buffer[154][6] ) );
  DFFQXL \row1_buffer_reg[153][6]  ( .D(\row1_buffer[154][6] ), .CK(clk), .Q(
        \row1_buffer[153][6] ) );
  DFFQXL \row1_buffer_reg[152][6]  ( .D(\row1_buffer[153][6] ), .CK(clk), .Q(
        \row1_buffer[152][6] ) );
  DFFQXL \row1_buffer_reg[151][6]  ( .D(\row1_buffer[152][6] ), .CK(clk), .Q(
        \row1_buffer[151][6] ) );
  DFFQXL \row1_buffer_reg[150][6]  ( .D(\row1_buffer[151][6] ), .CK(clk), .Q(
        \row1_buffer[150][6] ) );
  DFFQXL \row1_buffer_reg[149][6]  ( .D(\row1_buffer[150][6] ), .CK(clk), .Q(
        \row1_buffer[149][6] ) );
  DFFQXL \row1_buffer_reg[148][6]  ( .D(\row1_buffer[149][6] ), .CK(clk), .Q(
        \row1_buffer[148][6] ) );
  DFFQXL \row1_buffer_reg[147][6]  ( .D(\row1_buffer[148][6] ), .CK(clk), .Q(
        \row1_buffer[147][6] ) );
  DFFQXL \row1_buffer_reg[146][6]  ( .D(\row1_buffer[147][6] ), .CK(clk), .Q(
        \row1_buffer[146][6] ) );
  DFFQXL \row1_buffer_reg[145][6]  ( .D(\row1_buffer[146][6] ), .CK(clk), .Q(
        \row1_buffer[145][6] ) );
  DFFQXL \row1_buffer_reg[144][6]  ( .D(\row1_buffer[145][6] ), .CK(clk), .Q(
        \row1_buffer[144][6] ) );
  DFFQXL \row1_buffer_reg[143][6]  ( .D(\row1_buffer[144][6] ), .CK(clk), .Q(
        \row1_buffer[143][6] ) );
  DFFQXL \row1_buffer_reg[142][6]  ( .D(\row1_buffer[143][6] ), .CK(clk), .Q(
        \row1_buffer[142][6] ) );
  DFFQXL \row1_buffer_reg[141][6]  ( .D(\row1_buffer[142][6] ), .CK(clk), .Q(
        \row1_buffer[141][6] ) );
  DFFQXL \row1_buffer_reg[140][6]  ( .D(\row1_buffer[141][6] ), .CK(clk), .Q(
        \row1_buffer[140][6] ) );
  DFFQXL \row1_buffer_reg[139][6]  ( .D(\row1_buffer[140][6] ), .CK(clk), .Q(
        \row1_buffer[139][6] ) );
  DFFQXL \row1_buffer_reg[138][6]  ( .D(\row1_buffer[139][6] ), .CK(clk), .Q(
        \row1_buffer[138][6] ) );
  DFFQXL \row1_buffer_reg[137][6]  ( .D(\row1_buffer[138][6] ), .CK(clk), .Q(
        \row1_buffer[137][6] ) );
  DFFQXL \row1_buffer_reg[136][6]  ( .D(\row1_buffer[137][6] ), .CK(clk), .Q(
        \row1_buffer[136][6] ) );
  DFFQXL \row1_buffer_reg[135][6]  ( .D(\row1_buffer[136][6] ), .CK(clk), .Q(
        \row1_buffer[135][6] ) );
  DFFQXL \row1_buffer_reg[134][6]  ( .D(\row1_buffer[135][6] ), .CK(clk), .Q(
        \row1_buffer[134][6] ) );
  DFFQXL \row1_buffer_reg[133][6]  ( .D(\row1_buffer[134][6] ), .CK(clk), .Q(
        \row1_buffer[133][6] ) );
  DFFQXL \row1_buffer_reg[132][6]  ( .D(\row1_buffer[133][6] ), .CK(clk), .Q(
        \row1_buffer[132][6] ) );
  DFFQXL \row1_buffer_reg[131][6]  ( .D(\row1_buffer[132][6] ), .CK(clk), .Q(
        \row1_buffer[131][6] ) );
  DFFQXL \row1_buffer_reg[130][6]  ( .D(\row1_buffer[131][6] ), .CK(clk), .Q(
        \row1_buffer[130][6] ) );
  DFFQXL \row1_buffer_reg[129][6]  ( .D(\row1_buffer[130][6] ), .CK(clk), .Q(
        \row1_buffer[129][6] ) );
  DFFQXL \row1_buffer_reg[128][6]  ( .D(\row1_buffer[129][6] ), .CK(clk), .Q(
        \row1_buffer[128][6] ) );
  DFFQXL \row1_buffer_reg[127][6]  ( .D(\row1_buffer[128][6] ), .CK(clk), .Q(
        \row1_buffer[127][6] ) );
  DFFQXL \row1_buffer_reg[126][6]  ( .D(\row1_buffer[127][6] ), .CK(clk), .Q(
        \row1_buffer[126][6] ) );
  DFFQXL \row1_buffer_reg[125][6]  ( .D(\row1_buffer[126][6] ), .CK(clk), .Q(
        \row1_buffer[125][6] ) );
  DFFQXL \row1_buffer_reg[124][6]  ( .D(\row1_buffer[125][6] ), .CK(clk), .Q(
        \row1_buffer[124][6] ) );
  DFFQXL \row1_buffer_reg[123][6]  ( .D(\row1_buffer[124][6] ), .CK(clk), .Q(
        \row1_buffer[123][6] ) );
  DFFQXL \row1_buffer_reg[122][6]  ( .D(\row1_buffer[123][6] ), .CK(clk), .Q(
        \row1_buffer[122][6] ) );
  DFFQXL \row1_buffer_reg[121][6]  ( .D(\row1_buffer[122][6] ), .CK(clk), .Q(
        \row1_buffer[121][6] ) );
  DFFQXL \row1_buffer_reg[120][6]  ( .D(\row1_buffer[121][6] ), .CK(clk), .Q(
        \row1_buffer[120][6] ) );
  DFFQXL \row1_buffer_reg[119][6]  ( .D(\row1_buffer[120][6] ), .CK(clk), .Q(
        \row1_buffer[119][6] ) );
  DFFQXL \row1_buffer_reg[118][6]  ( .D(\row1_buffer[119][6] ), .CK(clk), .Q(
        \row1_buffer[118][6] ) );
  DFFQXL \row1_buffer_reg[117][6]  ( .D(\row1_buffer[118][6] ), .CK(clk), .Q(
        \row1_buffer[117][6] ) );
  DFFQXL \row1_buffer_reg[116][6]  ( .D(\row1_buffer[117][6] ), .CK(clk), .Q(
        \row1_buffer[116][6] ) );
  DFFQXL \row1_buffer_reg[115][6]  ( .D(\row1_buffer[116][6] ), .CK(clk), .Q(
        \row1_buffer[115][6] ) );
  DFFQXL \row1_buffer_reg[114][6]  ( .D(\row1_buffer[115][6] ), .CK(clk), .Q(
        \row1_buffer[114][6] ) );
  DFFQXL \row1_buffer_reg[113][6]  ( .D(\row1_buffer[114][6] ), .CK(clk), .Q(
        \row1_buffer[113][6] ) );
  DFFQXL \row1_buffer_reg[112][6]  ( .D(\row1_buffer[113][6] ), .CK(clk), .Q(
        \row1_buffer[112][6] ) );
  DFFQXL \row1_buffer_reg[111][6]  ( .D(\row1_buffer[112][6] ), .CK(clk), .Q(
        \row1_buffer[111][6] ) );
  DFFQXL \row1_buffer_reg[110][6]  ( .D(\row1_buffer[111][6] ), .CK(clk), .Q(
        \row1_buffer[110][6] ) );
  DFFQXL \row1_buffer_reg[109][6]  ( .D(\row1_buffer[110][6] ), .CK(clk), .Q(
        \row1_buffer[109][6] ) );
  DFFQXL \row1_buffer_reg[108][6]  ( .D(\row1_buffer[109][6] ), .CK(clk), .Q(
        \row1_buffer[108][6] ) );
  DFFQXL \row1_buffer_reg[107][6]  ( .D(\row1_buffer[108][6] ), .CK(clk), .Q(
        \row1_buffer[107][6] ) );
  DFFQXL \row1_buffer_reg[106][6]  ( .D(\row1_buffer[107][6] ), .CK(clk), .Q(
        \row1_buffer[106][6] ) );
  DFFQXL \row1_buffer_reg[105][6]  ( .D(\row1_buffer[106][6] ), .CK(clk), .Q(
        \row1_buffer[105][6] ) );
  DFFQXL \row1_buffer_reg[104][6]  ( .D(\row1_buffer[105][6] ), .CK(clk), .Q(
        \row1_buffer[104][6] ) );
  DFFQXL \row1_buffer_reg[103][6]  ( .D(\row1_buffer[104][6] ), .CK(clk), .Q(
        \row1_buffer[103][6] ) );
  DFFQXL \row1_buffer_reg[102][6]  ( .D(\row1_buffer[103][6] ), .CK(clk), .Q(
        \row1_buffer[102][6] ) );
  DFFQXL \row1_buffer_reg[101][6]  ( .D(\row1_buffer[102][6] ), .CK(clk), .Q(
        \row1_buffer[101][6] ) );
  DFFQXL \row1_buffer_reg[100][6]  ( .D(\row1_buffer[101][6] ), .CK(clk), .Q(
        \row1_buffer[100][6] ) );
  DFFQXL \row1_buffer_reg[99][6]  ( .D(\row1_buffer[100][6] ), .CK(clk), .Q(
        \row1_buffer[99][6] ) );
  DFFQXL \row1_buffer_reg[98][6]  ( .D(\row1_buffer[99][6] ), .CK(clk), .Q(
        \row1_buffer[98][6] ) );
  DFFQXL \row1_buffer_reg[97][6]  ( .D(\row1_buffer[98][6] ), .CK(clk), .Q(
        \row1_buffer[97][6] ) );
  DFFQXL \row1_buffer_reg[96][6]  ( .D(\row1_buffer[97][6] ), .CK(clk), .Q(
        \row1_buffer[96][6] ) );
  DFFQXL \row1_buffer_reg[95][6]  ( .D(\row1_buffer[96][6] ), .CK(clk), .Q(
        \row1_buffer[95][6] ) );
  DFFQXL \row1_buffer_reg[94][6]  ( .D(\row1_buffer[95][6] ), .CK(clk), .Q(
        \row1_buffer[94][6] ) );
  DFFQXL \row1_buffer_reg[93][6]  ( .D(\row1_buffer[94][6] ), .CK(clk), .Q(
        \row1_buffer[93][6] ) );
  DFFQXL \row1_buffer_reg[92][6]  ( .D(\row1_buffer[93][6] ), .CK(clk), .Q(
        \row1_buffer[92][6] ) );
  DFFQXL \row1_buffer_reg[91][6]  ( .D(\row1_buffer[92][6] ), .CK(clk), .Q(
        \row1_buffer[91][6] ) );
  DFFQXL \row1_buffer_reg[90][6]  ( .D(\row1_buffer[91][6] ), .CK(clk), .Q(
        \row1_buffer[90][6] ) );
  DFFQXL \row1_buffer_reg[89][6]  ( .D(\row1_buffer[90][6] ), .CK(clk), .Q(
        \row1_buffer[89][6] ) );
  DFFQXL \row1_buffer_reg[88][6]  ( .D(\row1_buffer[89][6] ), .CK(clk), .Q(
        \row1_buffer[88][6] ) );
  DFFQXL \row1_buffer_reg[87][6]  ( .D(\row1_buffer[88][6] ), .CK(clk), .Q(
        \row1_buffer[87][6] ) );
  DFFQXL \row1_buffer_reg[86][6]  ( .D(\row1_buffer[87][6] ), .CK(clk), .Q(
        \row1_buffer[86][6] ) );
  DFFQXL \row1_buffer_reg[85][6]  ( .D(\row1_buffer[86][6] ), .CK(clk), .Q(
        \row1_buffer[85][6] ) );
  DFFQXL \row1_buffer_reg[84][6]  ( .D(\row1_buffer[85][6] ), .CK(clk), .Q(
        \row1_buffer[84][6] ) );
  DFFQXL \row1_buffer_reg[83][6]  ( .D(\row1_buffer[84][6] ), .CK(clk), .Q(
        \row1_buffer[83][6] ) );
  DFFQXL \row1_buffer_reg[82][6]  ( .D(\row1_buffer[83][6] ), .CK(clk), .Q(
        \row1_buffer[82][6] ) );
  DFFQXL \row1_buffer_reg[81][6]  ( .D(\row1_buffer[82][6] ), .CK(clk), .Q(
        \row1_buffer[81][6] ) );
  DFFQXL \row1_buffer_reg[80][6]  ( .D(\row1_buffer[81][6] ), .CK(clk), .Q(
        \row1_buffer[80][6] ) );
  DFFQXL \row1_buffer_reg[79][6]  ( .D(\row1_buffer[80][6] ), .CK(clk), .Q(
        \row1_buffer[79][6] ) );
  DFFQXL \row1_buffer_reg[78][6]  ( .D(\row1_buffer[79][6] ), .CK(clk), .Q(
        \row1_buffer[78][6] ) );
  DFFQXL \row1_buffer_reg[77][6]  ( .D(\row1_buffer[78][6] ), .CK(clk), .Q(
        \row1_buffer[77][6] ) );
  DFFQXL \row1_buffer_reg[76][6]  ( .D(\row1_buffer[77][6] ), .CK(clk), .Q(
        \row1_buffer[76][6] ) );
  DFFQXL \row1_buffer_reg[75][6]  ( .D(\row1_buffer[76][6] ), .CK(clk), .Q(
        \row1_buffer[75][6] ) );
  DFFQXL \row1_buffer_reg[74][6]  ( .D(\row1_buffer[75][6] ), .CK(clk), .Q(
        \row1_buffer[74][6] ) );
  DFFQXL \row1_buffer_reg[73][6]  ( .D(\row1_buffer[74][6] ), .CK(clk), .Q(
        \row1_buffer[73][6] ) );
  DFFQXL \row1_buffer_reg[72][6]  ( .D(\row1_buffer[73][6] ), .CK(clk), .Q(
        \row1_buffer[72][6] ) );
  DFFQXL \row1_buffer_reg[71][6]  ( .D(\row1_buffer[72][6] ), .CK(clk), .Q(
        \row1_buffer[71][6] ) );
  DFFQXL \row1_buffer_reg[70][6]  ( .D(\row1_buffer[71][6] ), .CK(clk), .Q(
        \row1_buffer[70][6] ) );
  DFFQXL \row1_buffer_reg[69][6]  ( .D(\row1_buffer[70][6] ), .CK(clk), .Q(
        \row1_buffer[69][6] ) );
  DFFQXL \row1_buffer_reg[68][6]  ( .D(\row1_buffer[69][6] ), .CK(clk), .Q(
        \row1_buffer[68][6] ) );
  DFFQXL \row1_buffer_reg[67][6]  ( .D(\row1_buffer[68][6] ), .CK(clk), .Q(
        \row1_buffer[67][6] ) );
  DFFQXL \row1_buffer_reg[66][6]  ( .D(\row1_buffer[67][6] ), .CK(clk), .Q(
        \row1_buffer[66][6] ) );
  DFFQXL \row1_buffer_reg[65][6]  ( .D(\row1_buffer[66][6] ), .CK(clk), .Q(
        \row1_buffer[65][6] ) );
  DFFQXL \row1_buffer_reg[64][6]  ( .D(\row1_buffer[65][6] ), .CK(clk), .Q(
        \row1_buffer[64][6] ) );
  DFFQXL \row1_buffer_reg[63][6]  ( .D(\row1_buffer[64][6] ), .CK(clk), .Q(
        \row1_buffer[63][6] ) );
  DFFQXL \row1_buffer_reg[62][6]  ( .D(\row1_buffer[63][6] ), .CK(clk), .Q(
        \row1_buffer[62][6] ) );
  DFFQXL \row1_buffer_reg[61][6]  ( .D(\row1_buffer[62][6] ), .CK(clk), .Q(
        \row1_buffer[61][6] ) );
  DFFQXL \row1_buffer_reg[60][6]  ( .D(\row1_buffer[61][6] ), .CK(clk), .Q(
        \row1_buffer[60][6] ) );
  DFFQXL \row1_buffer_reg[59][6]  ( .D(\row1_buffer[60][6] ), .CK(clk), .Q(
        \row1_buffer[59][6] ) );
  DFFQXL \row1_buffer_reg[58][6]  ( .D(\row1_buffer[59][6] ), .CK(clk), .Q(
        \row1_buffer[58][6] ) );
  DFFQXL \row1_buffer_reg[57][6]  ( .D(\row1_buffer[58][6] ), .CK(clk), .Q(
        \row1_buffer[57][6] ) );
  DFFQXL \row1_buffer_reg[56][6]  ( .D(\row1_buffer[57][6] ), .CK(clk), .Q(
        \row1_buffer[56][6] ) );
  DFFQXL \row1_buffer_reg[55][6]  ( .D(\row1_buffer[56][6] ), .CK(clk), .Q(
        \row1_buffer[55][6] ) );
  DFFQXL \row1_buffer_reg[54][6]  ( .D(\row1_buffer[55][6] ), .CK(clk), .Q(
        \row1_buffer[54][6] ) );
  DFFQXL \row1_buffer_reg[53][6]  ( .D(\row1_buffer[54][6] ), .CK(clk), .Q(
        \row1_buffer[53][6] ) );
  DFFQXL \row1_buffer_reg[52][6]  ( .D(\row1_buffer[53][6] ), .CK(clk), .Q(
        \row1_buffer[52][6] ) );
  DFFQXL \row1_buffer_reg[51][6]  ( .D(\row1_buffer[52][6] ), .CK(clk), .Q(
        \row1_buffer[51][6] ) );
  DFFQXL \row1_buffer_reg[50][6]  ( .D(\row1_buffer[51][6] ), .CK(clk), .Q(
        \row1_buffer[50][6] ) );
  DFFQXL \row1_buffer_reg[49][6]  ( .D(\row1_buffer[50][6] ), .CK(clk), .Q(
        \row1_buffer[49][6] ) );
  DFFQXL \row1_buffer_reg[48][6]  ( .D(\row1_buffer[49][6] ), .CK(clk), .Q(
        \row1_buffer[48][6] ) );
  DFFQXL \row1_buffer_reg[47][6]  ( .D(\row1_buffer[48][6] ), .CK(clk), .Q(
        \row1_buffer[47][6] ) );
  DFFQXL \row1_buffer_reg[46][6]  ( .D(\row1_buffer[47][6] ), .CK(clk), .Q(
        \row1_buffer[46][6] ) );
  DFFQXL \row1_buffer_reg[45][6]  ( .D(\row1_buffer[46][6] ), .CK(clk), .Q(
        \row1_buffer[45][6] ) );
  DFFQXL \row1_buffer_reg[44][6]  ( .D(\row1_buffer[45][6] ), .CK(clk), .Q(
        \row1_buffer[44][6] ) );
  DFFQXL \row1_buffer_reg[43][6]  ( .D(\row1_buffer[44][6] ), .CK(clk), .Q(
        \row1_buffer[43][6] ) );
  DFFQXL \row1_buffer_reg[42][6]  ( .D(\row1_buffer[43][6] ), .CK(clk), .Q(
        \row1_buffer[42][6] ) );
  DFFQXL \row1_buffer_reg[41][6]  ( .D(\row1_buffer[42][6] ), .CK(clk), .Q(
        \row1_buffer[41][6] ) );
  DFFQXL \row1_buffer_reg[40][6]  ( .D(\row1_buffer[41][6] ), .CK(clk), .Q(
        \row1_buffer[40][6] ) );
  DFFQXL \row1_buffer_reg[39][6]  ( .D(\row1_buffer[40][6] ), .CK(clk), .Q(
        \row1_buffer[39][6] ) );
  DFFQXL \row1_buffer_reg[38][6]  ( .D(\row1_buffer[39][6] ), .CK(clk), .Q(
        \row1_buffer[38][6] ) );
  DFFQXL \row1_buffer_reg[37][6]  ( .D(\row1_buffer[38][6] ), .CK(clk), .Q(
        \row1_buffer[37][6] ) );
  DFFQXL \row1_buffer_reg[36][6]  ( .D(\row1_buffer[37][6] ), .CK(clk), .Q(
        \row1_buffer[36][6] ) );
  DFFQXL \row1_buffer_reg[35][6]  ( .D(\row1_buffer[36][6] ), .CK(clk), .Q(
        \row1_buffer[35][6] ) );
  DFFQXL \row1_buffer_reg[34][6]  ( .D(\row1_buffer[35][6] ), .CK(clk), .Q(
        \row1_buffer[34][6] ) );
  DFFQXL \row1_buffer_reg[33][6]  ( .D(\row1_buffer[34][6] ), .CK(clk), .Q(
        \row1_buffer[33][6] ) );
  DFFQXL \row1_buffer_reg[32][6]  ( .D(\row1_buffer[33][6] ), .CK(clk), .Q(
        \row1_buffer[32][6] ) );
  DFFQXL \row1_buffer_reg[31][6]  ( .D(\row1_buffer[32][6] ), .CK(clk), .Q(
        \row1_buffer[31][6] ) );
  DFFQXL \row1_buffer_reg[30][6]  ( .D(\row1_buffer[31][6] ), .CK(clk), .Q(
        \row1_buffer[30][6] ) );
  DFFQXL \row1_buffer_reg[29][6]  ( .D(\row1_buffer[30][6] ), .CK(clk), .Q(
        \row1_buffer[29][6] ) );
  DFFQXL \row1_buffer_reg[28][6]  ( .D(\row1_buffer[29][6] ), .CK(clk), .Q(
        \row1_buffer[28][6] ) );
  DFFQXL \row1_buffer_reg[27][6]  ( .D(\row1_buffer[28][6] ), .CK(clk), .Q(
        \row1_buffer[27][6] ) );
  DFFQXL \row1_buffer_reg[26][6]  ( .D(\row1_buffer[27][6] ), .CK(clk), .Q(
        \row1_buffer[26][6] ) );
  DFFQXL \row1_buffer_reg[25][6]  ( .D(\row1_buffer[26][6] ), .CK(clk), .Q(
        \row1_buffer[25][6] ) );
  DFFQXL \row1_buffer_reg[24][6]  ( .D(\row1_buffer[25][6] ), .CK(clk), .Q(
        \row1_buffer[24][6] ) );
  DFFQXL \row1_buffer_reg[23][6]  ( .D(\row1_buffer[24][6] ), .CK(clk), .Q(
        \row1_buffer[23][6] ) );
  DFFQXL \row1_buffer_reg[22][6]  ( .D(\row1_buffer[23][6] ), .CK(clk), .Q(
        \row1_buffer[22][6] ) );
  DFFQXL \row1_buffer_reg[21][6]  ( .D(\row1_buffer[22][6] ), .CK(clk), .Q(
        \row1_buffer[21][6] ) );
  DFFQXL \row1_buffer_reg[20][6]  ( .D(\row1_buffer[21][6] ), .CK(clk), .Q(
        \row1_buffer[20][6] ) );
  DFFQXL \row1_buffer_reg[19][6]  ( .D(\row1_buffer[20][6] ), .CK(clk), .Q(
        \row1_buffer[19][6] ) );
  DFFQXL \row1_buffer_reg[18][6]  ( .D(\row1_buffer[19][6] ), .CK(clk), .Q(
        \row1_buffer[18][6] ) );
  DFFQXL \row1_buffer_reg[17][6]  ( .D(\row1_buffer[18][6] ), .CK(clk), .Q(
        \row1_buffer[17][6] ) );
  DFFQXL \row1_buffer_reg[16][6]  ( .D(\row1_buffer[17][6] ), .CK(clk), .Q(
        \row1_buffer[16][6] ) );
  DFFQXL \row1_buffer_reg[15][6]  ( .D(\row1_buffer[16][6] ), .CK(clk), .Q(
        \row1_buffer[15][6] ) );
  DFFQXL \row1_buffer_reg[14][6]  ( .D(\row1_buffer[15][6] ), .CK(clk), .Q(
        \row1_buffer[14][6] ) );
  DFFQXL \row1_buffer_reg[13][6]  ( .D(\row1_buffer[14][6] ), .CK(clk), .Q(
        \row1_buffer[13][6] ) );
  DFFQXL \row1_buffer_reg[12][6]  ( .D(\row1_buffer[13][6] ), .CK(clk), .Q(
        \row1_buffer[12][6] ) );
  DFFQXL \row1_buffer_reg[11][6]  ( .D(\row1_buffer[12][6] ), .CK(clk), .Q(
        \row1_buffer[11][6] ) );
  DFFQXL \row1_buffer_reg[10][6]  ( .D(\row1_buffer[11][6] ), .CK(clk), .Q(
        \row1_buffer[10][6] ) );
  DFFQXL \row1_buffer_reg[9][6]  ( .D(\row1_buffer[10][6] ), .CK(clk), .Q(
        \row1_buffer[9][6] ) );
  DFFQXL \row1_buffer_reg[8][6]  ( .D(\row1_buffer[9][6] ), .CK(clk), .Q(
        \row1_buffer[8][6] ) );
  DFFQXL \row1_buffer_reg[7][6]  ( .D(\row1_buffer[8][6] ), .CK(clk), .Q(
        \row1_buffer[7][6] ) );
  DFFQXL \row1_buffer_reg[6][6]  ( .D(\row1_buffer[7][6] ), .CK(clk), .Q(
        \row1_buffer[6][6] ) );
  DFFQXL \row1_buffer_reg[5][6]  ( .D(\row1_buffer[6][6] ), .CK(clk), .Q(
        \row1_buffer[5][6] ) );
  DFFQXL \row1_buffer_reg[4][6]  ( .D(\row1_buffer[5][6] ), .CK(clk), .Q(
        \row1_buffer[4][6] ) );
  DFFQXL \row1_buffer_reg[3][6]  ( .D(\row1_buffer[4][6] ), .CK(clk), .Q(
        \row1_buffer[3][6] ) );
  DFFQXL \row2_buffer_reg[225][5]  ( .D(\row3_buffer[0][5] ), .CK(clk), .Q(
        \row2_buffer[225][5] ) );
  DFFQXL \row2_buffer_reg[224][5]  ( .D(\row2_buffer[225][5] ), .CK(clk), .Q(
        \row2_buffer[224][5] ) );
  DFFQXL \row2_buffer_reg[223][5]  ( .D(\row2_buffer[224][5] ), .CK(clk), .Q(
        \row2_buffer[223][5] ) );
  DFFQXL \row2_buffer_reg[222][5]  ( .D(\row2_buffer[223][5] ), .CK(clk), .Q(
        \row2_buffer[222][5] ) );
  DFFQXL \row2_buffer_reg[221][5]  ( .D(\row2_buffer[222][5] ), .CK(clk), .Q(
        \row2_buffer[221][5] ) );
  DFFQXL \row2_buffer_reg[220][5]  ( .D(\row2_buffer[221][5] ), .CK(clk), .Q(
        \row2_buffer[220][5] ) );
  DFFQXL \row2_buffer_reg[219][5]  ( .D(\row2_buffer[220][5] ), .CK(clk), .Q(
        \row2_buffer[219][5] ) );
  DFFQXL \row2_buffer_reg[218][5]  ( .D(\row2_buffer[219][5] ), .CK(clk), .Q(
        \row2_buffer[218][5] ) );
  DFFQXL \row2_buffer_reg[217][5]  ( .D(\row2_buffer[218][5] ), .CK(clk), .Q(
        \row2_buffer[217][5] ) );
  DFFQXL \row2_buffer_reg[216][5]  ( .D(\row2_buffer[217][5] ), .CK(clk), .Q(
        \row2_buffer[216][5] ) );
  DFFQXL \row2_buffer_reg[215][5]  ( .D(\row2_buffer[216][5] ), .CK(clk), .Q(
        \row2_buffer[215][5] ) );
  DFFQXL \row2_buffer_reg[214][5]  ( .D(\row2_buffer[215][5] ), .CK(clk), .Q(
        \row2_buffer[214][5] ) );
  DFFQXL \row2_buffer_reg[213][5]  ( .D(\row2_buffer[214][5] ), .CK(clk), .Q(
        \row2_buffer[213][5] ) );
  DFFQXL \row2_buffer_reg[212][5]  ( .D(\row2_buffer[213][5] ), .CK(clk), .Q(
        \row2_buffer[212][5] ) );
  DFFQXL \row2_buffer_reg[211][5]  ( .D(\row2_buffer[212][5] ), .CK(clk), .Q(
        \row2_buffer[211][5] ) );
  DFFQXL \row2_buffer_reg[210][5]  ( .D(\row2_buffer[211][5] ), .CK(clk), .Q(
        \row2_buffer[210][5] ) );
  DFFQXL \row2_buffer_reg[209][5]  ( .D(\row2_buffer[210][5] ), .CK(clk), .Q(
        \row2_buffer[209][5] ) );
  DFFQXL \row2_buffer_reg[208][5]  ( .D(\row2_buffer[209][5] ), .CK(clk), .Q(
        \row2_buffer[208][5] ) );
  DFFQXL \row2_buffer_reg[207][5]  ( .D(\row2_buffer[208][5] ), .CK(clk), .Q(
        \row2_buffer[207][5] ) );
  DFFQXL \row2_buffer_reg[206][5]  ( .D(\row2_buffer[207][5] ), .CK(clk), .Q(
        \row2_buffer[206][5] ) );
  DFFQXL \row2_buffer_reg[205][5]  ( .D(\row2_buffer[206][5] ), .CK(clk), .Q(
        \row2_buffer[205][5] ) );
  DFFQXL \row2_buffer_reg[204][5]  ( .D(\row2_buffer[205][5] ), .CK(clk), .Q(
        \row2_buffer[204][5] ) );
  DFFQXL \row2_buffer_reg[203][5]  ( .D(\row2_buffer[204][5] ), .CK(clk), .Q(
        \row2_buffer[203][5] ) );
  DFFQXL \row2_buffer_reg[202][5]  ( .D(\row2_buffer[203][5] ), .CK(clk), .Q(
        \row2_buffer[202][5] ) );
  DFFQXL \row2_buffer_reg[201][5]  ( .D(\row2_buffer[202][5] ), .CK(clk), .Q(
        \row2_buffer[201][5] ) );
  DFFQXL \row2_buffer_reg[200][5]  ( .D(\row2_buffer[201][5] ), .CK(clk), .Q(
        \row2_buffer[200][5] ) );
  DFFQXL \row2_buffer_reg[199][5]  ( .D(\row2_buffer[200][5] ), .CK(clk), .Q(
        \row2_buffer[199][5] ) );
  DFFQXL \row2_buffer_reg[198][5]  ( .D(\row2_buffer[199][5] ), .CK(clk), .Q(
        \row2_buffer[198][5] ) );
  DFFQXL \row2_buffer_reg[197][5]  ( .D(\row2_buffer[198][5] ), .CK(clk), .Q(
        \row2_buffer[197][5] ) );
  DFFQXL \row2_buffer_reg[196][5]  ( .D(\row2_buffer[197][5] ), .CK(clk), .Q(
        \row2_buffer[196][5] ) );
  DFFQXL \row2_buffer_reg[195][5]  ( .D(\row2_buffer[196][5] ), .CK(clk), .Q(
        \row2_buffer[195][5] ) );
  DFFQXL \row2_buffer_reg[194][5]  ( .D(\row2_buffer[195][5] ), .CK(clk), .Q(
        \row2_buffer[194][5] ) );
  DFFQXL \row2_buffer_reg[193][5]  ( .D(\row2_buffer[194][5] ), .CK(clk), .Q(
        \row2_buffer[193][5] ) );
  DFFQXL \row2_buffer_reg[192][5]  ( .D(\row2_buffer[193][5] ), .CK(clk), .Q(
        \row2_buffer[192][5] ) );
  DFFQXL \row2_buffer_reg[191][5]  ( .D(\row2_buffer[192][5] ), .CK(clk), .Q(
        \row2_buffer[191][5] ) );
  DFFQXL \row2_buffer_reg[190][5]  ( .D(\row2_buffer[191][5] ), .CK(clk), .Q(
        \row2_buffer[190][5] ) );
  DFFQXL \row2_buffer_reg[189][5]  ( .D(\row2_buffer[190][5] ), .CK(clk), .Q(
        \row2_buffer[189][5] ) );
  DFFQXL \row2_buffer_reg[188][5]  ( .D(\row2_buffer[189][5] ), .CK(clk), .Q(
        \row2_buffer[188][5] ) );
  DFFQXL \row2_buffer_reg[187][5]  ( .D(\row2_buffer[188][5] ), .CK(clk), .Q(
        \row2_buffer[187][5] ) );
  DFFQXL \row2_buffer_reg[186][5]  ( .D(\row2_buffer[187][5] ), .CK(clk), .Q(
        \row2_buffer[186][5] ) );
  DFFQXL \row2_buffer_reg[185][5]  ( .D(\row2_buffer[186][5] ), .CK(clk), .Q(
        \row2_buffer[185][5] ) );
  DFFQXL \row2_buffer_reg[184][5]  ( .D(\row2_buffer[185][5] ), .CK(clk), .Q(
        \row2_buffer[184][5] ) );
  DFFQXL \row2_buffer_reg[183][5]  ( .D(\row2_buffer[184][5] ), .CK(clk), .Q(
        \row2_buffer[183][5] ) );
  DFFQXL \row2_buffer_reg[182][5]  ( .D(\row2_buffer[183][5] ), .CK(clk), .Q(
        \row2_buffer[182][5] ) );
  DFFQXL \row2_buffer_reg[181][5]  ( .D(\row2_buffer[182][5] ), .CK(clk), .Q(
        \row2_buffer[181][5] ) );
  DFFQXL \row2_buffer_reg[180][5]  ( .D(\row2_buffer[181][5] ), .CK(clk), .Q(
        \row2_buffer[180][5] ) );
  DFFQXL \row2_buffer_reg[179][5]  ( .D(\row2_buffer[180][5] ), .CK(clk), .Q(
        \row2_buffer[179][5] ) );
  DFFQXL \row2_buffer_reg[178][5]  ( .D(\row2_buffer[179][5] ), .CK(clk), .Q(
        \row2_buffer[178][5] ) );
  DFFQXL \row2_buffer_reg[177][5]  ( .D(\row2_buffer[178][5] ), .CK(clk), .Q(
        \row2_buffer[177][5] ) );
  DFFQXL \row2_buffer_reg[176][5]  ( .D(\row2_buffer[177][5] ), .CK(clk), .Q(
        \row2_buffer[176][5] ) );
  DFFQXL \row2_buffer_reg[175][5]  ( .D(\row2_buffer[176][5] ), .CK(clk), .Q(
        \row2_buffer[175][5] ) );
  DFFQXL \row2_buffer_reg[174][5]  ( .D(\row2_buffer[175][5] ), .CK(clk), .Q(
        \row2_buffer[174][5] ) );
  DFFQXL \row2_buffer_reg[173][5]  ( .D(\row2_buffer[174][5] ), .CK(clk), .Q(
        \row2_buffer[173][5] ) );
  DFFQXL \row2_buffer_reg[172][5]  ( .D(\row2_buffer[173][5] ), .CK(clk), .Q(
        \row2_buffer[172][5] ) );
  DFFQXL \row2_buffer_reg[171][5]  ( .D(\row2_buffer[172][5] ), .CK(clk), .Q(
        \row2_buffer[171][5] ) );
  DFFQXL \row2_buffer_reg[170][5]  ( .D(\row2_buffer[171][5] ), .CK(clk), .Q(
        \row2_buffer[170][5] ) );
  DFFQXL \row2_buffer_reg[169][5]  ( .D(\row2_buffer[170][5] ), .CK(clk), .Q(
        \row2_buffer[169][5] ) );
  DFFQXL \row2_buffer_reg[168][5]  ( .D(\row2_buffer[169][5] ), .CK(clk), .Q(
        \row2_buffer[168][5] ) );
  DFFQXL \row2_buffer_reg[167][5]  ( .D(\row2_buffer[168][5] ), .CK(clk), .Q(
        \row2_buffer[167][5] ) );
  DFFQXL \row2_buffer_reg[166][5]  ( .D(\row2_buffer[167][5] ), .CK(clk), .Q(
        \row2_buffer[166][5] ) );
  DFFQXL \row2_buffer_reg[165][5]  ( .D(\row2_buffer[166][5] ), .CK(clk), .Q(
        \row2_buffer[165][5] ) );
  DFFQXL \row2_buffer_reg[164][5]  ( .D(\row2_buffer[165][5] ), .CK(clk), .Q(
        \row2_buffer[164][5] ) );
  DFFQXL \row2_buffer_reg[163][5]  ( .D(\row2_buffer[164][5] ), .CK(clk), .Q(
        \row2_buffer[163][5] ) );
  DFFQXL \row2_buffer_reg[162][5]  ( .D(\row2_buffer[163][5] ), .CK(clk), .Q(
        \row2_buffer[162][5] ) );
  DFFQXL \row2_buffer_reg[161][5]  ( .D(\row2_buffer[162][5] ), .CK(clk), .Q(
        \row2_buffer[161][5] ) );
  DFFQXL \row2_buffer_reg[160][5]  ( .D(\row2_buffer[161][5] ), .CK(clk), .Q(
        \row2_buffer[160][5] ) );
  DFFQXL \row2_buffer_reg[159][5]  ( .D(\row2_buffer[160][5] ), .CK(clk), .Q(
        \row2_buffer[159][5] ) );
  DFFQXL \row2_buffer_reg[158][5]  ( .D(\row2_buffer[159][5] ), .CK(clk), .Q(
        \row2_buffer[158][5] ) );
  DFFQXL \row2_buffer_reg[157][5]  ( .D(\row2_buffer[158][5] ), .CK(clk), .Q(
        \row2_buffer[157][5] ) );
  DFFQXL \row2_buffer_reg[156][5]  ( .D(\row2_buffer[157][5] ), .CK(clk), .Q(
        \row2_buffer[156][5] ) );
  DFFQXL \row2_buffer_reg[155][5]  ( .D(\row2_buffer[156][5] ), .CK(clk), .Q(
        \row2_buffer[155][5] ) );
  DFFQXL \row2_buffer_reg[154][5]  ( .D(\row2_buffer[155][5] ), .CK(clk), .Q(
        \row2_buffer[154][5] ) );
  DFFQXL \row2_buffer_reg[153][5]  ( .D(\row2_buffer[154][5] ), .CK(clk), .Q(
        \row2_buffer[153][5] ) );
  DFFQXL \row2_buffer_reg[152][5]  ( .D(\row2_buffer[153][5] ), .CK(clk), .Q(
        \row2_buffer[152][5] ) );
  DFFQXL \row2_buffer_reg[151][5]  ( .D(\row2_buffer[152][5] ), .CK(clk), .Q(
        \row2_buffer[151][5] ) );
  DFFQXL \row2_buffer_reg[150][5]  ( .D(\row2_buffer[151][5] ), .CK(clk), .Q(
        \row2_buffer[150][5] ) );
  DFFQXL \row2_buffer_reg[149][5]  ( .D(\row2_buffer[150][5] ), .CK(clk), .Q(
        \row2_buffer[149][5] ) );
  DFFQXL \row2_buffer_reg[148][5]  ( .D(\row2_buffer[149][5] ), .CK(clk), .Q(
        \row2_buffer[148][5] ) );
  DFFQXL \row2_buffer_reg[147][5]  ( .D(\row2_buffer[148][5] ), .CK(clk), .Q(
        \row2_buffer[147][5] ) );
  DFFQXL \row2_buffer_reg[146][5]  ( .D(\row2_buffer[147][5] ), .CK(clk), .Q(
        \row2_buffer[146][5] ) );
  DFFQXL \row2_buffer_reg[145][5]  ( .D(\row2_buffer[146][5] ), .CK(clk), .Q(
        \row2_buffer[145][5] ) );
  DFFQXL \row2_buffer_reg[144][5]  ( .D(\row2_buffer[145][5] ), .CK(clk), .Q(
        \row2_buffer[144][5] ) );
  DFFQXL \row2_buffer_reg[143][5]  ( .D(\row2_buffer[144][5] ), .CK(clk), .Q(
        \row2_buffer[143][5] ) );
  DFFQXL \row2_buffer_reg[142][5]  ( .D(\row2_buffer[143][5] ), .CK(clk), .Q(
        \row2_buffer[142][5] ) );
  DFFQXL \row2_buffer_reg[141][5]  ( .D(\row2_buffer[142][5] ), .CK(clk), .Q(
        \row2_buffer[141][5] ) );
  DFFQXL \row2_buffer_reg[140][5]  ( .D(\row2_buffer[141][5] ), .CK(clk), .Q(
        \row2_buffer[140][5] ) );
  DFFQXL \row2_buffer_reg[139][5]  ( .D(\row2_buffer[140][5] ), .CK(clk), .Q(
        \row2_buffer[139][5] ) );
  DFFQXL \row2_buffer_reg[138][5]  ( .D(\row2_buffer[139][5] ), .CK(clk), .Q(
        \row2_buffer[138][5] ) );
  DFFQXL \row2_buffer_reg[137][5]  ( .D(\row2_buffer[138][5] ), .CK(clk), .Q(
        \row2_buffer[137][5] ) );
  DFFQXL \row2_buffer_reg[136][5]  ( .D(\row2_buffer[137][5] ), .CK(clk), .Q(
        \row2_buffer[136][5] ) );
  DFFQXL \row2_buffer_reg[135][5]  ( .D(\row2_buffer[136][5] ), .CK(clk), .Q(
        \row2_buffer[135][5] ) );
  DFFQXL \row2_buffer_reg[134][5]  ( .D(\row2_buffer[135][5] ), .CK(clk), .Q(
        \row2_buffer[134][5] ) );
  DFFQXL \row2_buffer_reg[133][5]  ( .D(\row2_buffer[134][5] ), .CK(clk), .Q(
        \row2_buffer[133][5] ) );
  DFFQXL \row2_buffer_reg[132][5]  ( .D(\row2_buffer[133][5] ), .CK(clk), .Q(
        \row2_buffer[132][5] ) );
  DFFQXL \row2_buffer_reg[131][5]  ( .D(\row2_buffer[132][5] ), .CK(clk), .Q(
        \row2_buffer[131][5] ) );
  DFFQXL \row2_buffer_reg[130][5]  ( .D(\row2_buffer[131][5] ), .CK(clk), .Q(
        \row2_buffer[130][5] ) );
  DFFQXL \row2_buffer_reg[129][5]  ( .D(\row2_buffer[130][5] ), .CK(clk), .Q(
        \row2_buffer[129][5] ) );
  DFFQXL \row2_buffer_reg[128][5]  ( .D(\row2_buffer[129][5] ), .CK(clk), .Q(
        \row2_buffer[128][5] ) );
  DFFQXL \row2_buffer_reg[127][5]  ( .D(\row2_buffer[128][5] ), .CK(clk), .Q(
        \row2_buffer[127][5] ) );
  DFFQXL \row2_buffer_reg[126][5]  ( .D(\row2_buffer[127][5] ), .CK(clk), .Q(
        \row2_buffer[126][5] ) );
  DFFQXL \row2_buffer_reg[125][5]  ( .D(\row2_buffer[126][5] ), .CK(clk), .Q(
        \row2_buffer[125][5] ) );
  DFFQXL \row2_buffer_reg[124][5]  ( .D(\row2_buffer[125][5] ), .CK(clk), .Q(
        \row2_buffer[124][5] ) );
  DFFQXL \row2_buffer_reg[123][5]  ( .D(\row2_buffer[124][5] ), .CK(clk), .Q(
        \row2_buffer[123][5] ) );
  DFFQXL \row2_buffer_reg[122][5]  ( .D(\row2_buffer[123][5] ), .CK(clk), .Q(
        \row2_buffer[122][5] ) );
  DFFQXL \row2_buffer_reg[121][5]  ( .D(\row2_buffer[122][5] ), .CK(clk), .Q(
        \row2_buffer[121][5] ) );
  DFFQXL \row2_buffer_reg[120][5]  ( .D(\row2_buffer[121][5] ), .CK(clk), .Q(
        \row2_buffer[120][5] ) );
  DFFQXL \row2_buffer_reg[119][5]  ( .D(\row2_buffer[120][5] ), .CK(clk), .Q(
        \row2_buffer[119][5] ) );
  DFFQXL \row2_buffer_reg[118][5]  ( .D(\row2_buffer[119][5] ), .CK(clk), .Q(
        \row2_buffer[118][5] ) );
  DFFQXL \row2_buffer_reg[117][5]  ( .D(\row2_buffer[118][5] ), .CK(clk), .Q(
        \row2_buffer[117][5] ) );
  DFFQXL \row2_buffer_reg[116][5]  ( .D(\row2_buffer[117][5] ), .CK(clk), .Q(
        \row2_buffer[116][5] ) );
  DFFQXL \row2_buffer_reg[115][5]  ( .D(\row2_buffer[116][5] ), .CK(clk), .Q(
        \row2_buffer[115][5] ) );
  DFFQXL \row2_buffer_reg[114][5]  ( .D(\row2_buffer[115][5] ), .CK(clk), .Q(
        \row2_buffer[114][5] ) );
  DFFQXL \row2_buffer_reg[113][5]  ( .D(\row2_buffer[114][5] ), .CK(clk), .Q(
        \row2_buffer[113][5] ) );
  DFFQXL \row2_buffer_reg[112][5]  ( .D(\row2_buffer[113][5] ), .CK(clk), .Q(
        \row2_buffer[112][5] ) );
  DFFQXL \row2_buffer_reg[111][5]  ( .D(\row2_buffer[112][5] ), .CK(clk), .Q(
        \row2_buffer[111][5] ) );
  DFFQXL \row2_buffer_reg[110][5]  ( .D(\row2_buffer[111][5] ), .CK(clk), .Q(
        \row2_buffer[110][5] ) );
  DFFQXL \row2_buffer_reg[109][5]  ( .D(\row2_buffer[110][5] ), .CK(clk), .Q(
        \row2_buffer[109][5] ) );
  DFFQXL \row2_buffer_reg[108][5]  ( .D(\row2_buffer[109][5] ), .CK(clk), .Q(
        \row2_buffer[108][5] ) );
  DFFQXL \row2_buffer_reg[107][5]  ( .D(\row2_buffer[108][5] ), .CK(clk), .Q(
        \row2_buffer[107][5] ) );
  DFFQXL \row2_buffer_reg[106][5]  ( .D(\row2_buffer[107][5] ), .CK(clk), .Q(
        \row2_buffer[106][5] ) );
  DFFQXL \row2_buffer_reg[105][5]  ( .D(\row2_buffer[106][5] ), .CK(clk), .Q(
        \row2_buffer[105][5] ) );
  DFFQXL \row2_buffer_reg[104][5]  ( .D(\row2_buffer[105][5] ), .CK(clk), .Q(
        \row2_buffer[104][5] ) );
  DFFQXL \row2_buffer_reg[103][5]  ( .D(\row2_buffer[104][5] ), .CK(clk), .Q(
        \row2_buffer[103][5] ) );
  DFFQXL \row2_buffer_reg[102][5]  ( .D(\row2_buffer[103][5] ), .CK(clk), .Q(
        \row2_buffer[102][5] ) );
  DFFQXL \row2_buffer_reg[101][5]  ( .D(\row2_buffer[102][5] ), .CK(clk), .Q(
        \row2_buffer[101][5] ) );
  DFFQXL \row2_buffer_reg[100][5]  ( .D(\row2_buffer[101][5] ), .CK(clk), .Q(
        \row2_buffer[100][5] ) );
  DFFQXL \row2_buffer_reg[99][5]  ( .D(\row2_buffer[100][5] ), .CK(clk), .Q(
        \row2_buffer[99][5] ) );
  DFFQXL \row2_buffer_reg[98][5]  ( .D(\row2_buffer[99][5] ), .CK(clk), .Q(
        \row2_buffer[98][5] ) );
  DFFQXL \row2_buffer_reg[97][5]  ( .D(\row2_buffer[98][5] ), .CK(clk), .Q(
        \row2_buffer[97][5] ) );
  DFFQXL \row2_buffer_reg[96][5]  ( .D(\row2_buffer[97][5] ), .CK(clk), .Q(
        \row2_buffer[96][5] ) );
  DFFQXL \row2_buffer_reg[95][5]  ( .D(\row2_buffer[96][5] ), .CK(clk), .Q(
        \row2_buffer[95][5] ) );
  DFFQXL \row2_buffer_reg[94][5]  ( .D(\row2_buffer[95][5] ), .CK(clk), .Q(
        \row2_buffer[94][5] ) );
  DFFQXL \row2_buffer_reg[93][5]  ( .D(\row2_buffer[94][5] ), .CK(clk), .Q(
        \row2_buffer[93][5] ) );
  DFFQXL \row2_buffer_reg[92][5]  ( .D(\row2_buffer[93][5] ), .CK(clk), .Q(
        \row2_buffer[92][5] ) );
  DFFQXL \row2_buffer_reg[91][5]  ( .D(\row2_buffer[92][5] ), .CK(clk), .Q(
        \row2_buffer[91][5] ) );
  DFFQXL \row2_buffer_reg[90][5]  ( .D(\row2_buffer[91][5] ), .CK(clk), .Q(
        \row2_buffer[90][5] ) );
  DFFQXL \row2_buffer_reg[89][5]  ( .D(\row2_buffer[90][5] ), .CK(clk), .Q(
        \row2_buffer[89][5] ) );
  DFFQXL \row2_buffer_reg[88][5]  ( .D(\row2_buffer[89][5] ), .CK(clk), .Q(
        \row2_buffer[88][5] ) );
  DFFQXL \row2_buffer_reg[87][5]  ( .D(\row2_buffer[88][5] ), .CK(clk), .Q(
        \row2_buffer[87][5] ) );
  DFFQXL \row2_buffer_reg[86][5]  ( .D(\row2_buffer[87][5] ), .CK(clk), .Q(
        \row2_buffer[86][5] ) );
  DFFQXL \row2_buffer_reg[85][5]  ( .D(\row2_buffer[86][5] ), .CK(clk), .Q(
        \row2_buffer[85][5] ) );
  DFFQXL \row2_buffer_reg[84][5]  ( .D(\row2_buffer[85][5] ), .CK(clk), .Q(
        \row2_buffer[84][5] ) );
  DFFQXL \row2_buffer_reg[83][5]  ( .D(\row2_buffer[84][5] ), .CK(clk), .Q(
        \row2_buffer[83][5] ) );
  DFFQXL \row2_buffer_reg[82][5]  ( .D(\row2_buffer[83][5] ), .CK(clk), .Q(
        \row2_buffer[82][5] ) );
  DFFQXL \row2_buffer_reg[81][5]  ( .D(\row2_buffer[82][5] ), .CK(clk), .Q(
        \row2_buffer[81][5] ) );
  DFFQXL \row2_buffer_reg[80][5]  ( .D(\row2_buffer[81][5] ), .CK(clk), .Q(
        \row2_buffer[80][5] ) );
  DFFQXL \row2_buffer_reg[79][5]  ( .D(\row2_buffer[80][5] ), .CK(clk), .Q(
        \row2_buffer[79][5] ) );
  DFFQXL \row2_buffer_reg[78][5]  ( .D(\row2_buffer[79][5] ), .CK(clk), .Q(
        \row2_buffer[78][5] ) );
  DFFQXL \row2_buffer_reg[77][5]  ( .D(\row2_buffer[78][5] ), .CK(clk), .Q(
        \row2_buffer[77][5] ) );
  DFFQXL \row2_buffer_reg[76][5]  ( .D(\row2_buffer[77][5] ), .CK(clk), .Q(
        \row2_buffer[76][5] ) );
  DFFQXL \row2_buffer_reg[75][5]  ( .D(\row2_buffer[76][5] ), .CK(clk), .Q(
        \row2_buffer[75][5] ) );
  DFFQXL \row2_buffer_reg[74][5]  ( .D(\row2_buffer[75][5] ), .CK(clk), .Q(
        \row2_buffer[74][5] ) );
  DFFQXL \row2_buffer_reg[73][5]  ( .D(\row2_buffer[74][5] ), .CK(clk), .Q(
        \row2_buffer[73][5] ) );
  DFFQXL \row2_buffer_reg[72][5]  ( .D(\row2_buffer[73][5] ), .CK(clk), .Q(
        \row2_buffer[72][5] ) );
  DFFQXL \row2_buffer_reg[71][5]  ( .D(\row2_buffer[72][5] ), .CK(clk), .Q(
        \row2_buffer[71][5] ) );
  DFFQXL \row2_buffer_reg[70][5]  ( .D(\row2_buffer[71][5] ), .CK(clk), .Q(
        \row2_buffer[70][5] ) );
  DFFQXL \row2_buffer_reg[69][5]  ( .D(\row2_buffer[70][5] ), .CK(clk), .Q(
        \row2_buffer[69][5] ) );
  DFFQXL \row2_buffer_reg[68][5]  ( .D(\row2_buffer[69][5] ), .CK(clk), .Q(
        \row2_buffer[68][5] ) );
  DFFQXL \row2_buffer_reg[67][5]  ( .D(\row2_buffer[68][5] ), .CK(clk), .Q(
        \row2_buffer[67][5] ) );
  DFFQXL \row2_buffer_reg[66][5]  ( .D(\row2_buffer[67][5] ), .CK(clk), .Q(
        \row2_buffer[66][5] ) );
  DFFQXL \row2_buffer_reg[65][5]  ( .D(\row2_buffer[66][5] ), .CK(clk), .Q(
        \row2_buffer[65][5] ) );
  DFFQXL \row2_buffer_reg[64][5]  ( .D(\row2_buffer[65][5] ), .CK(clk), .Q(
        \row2_buffer[64][5] ) );
  DFFQXL \row2_buffer_reg[63][5]  ( .D(\row2_buffer[64][5] ), .CK(clk), .Q(
        \row2_buffer[63][5] ) );
  DFFQXL \row2_buffer_reg[62][5]  ( .D(\row2_buffer[63][5] ), .CK(clk), .Q(
        \row2_buffer[62][5] ) );
  DFFQXL \row2_buffer_reg[61][5]  ( .D(\row2_buffer[62][5] ), .CK(clk), .Q(
        \row2_buffer[61][5] ) );
  DFFQXL \row2_buffer_reg[60][5]  ( .D(\row2_buffer[61][5] ), .CK(clk), .Q(
        \row2_buffer[60][5] ) );
  DFFQXL \row2_buffer_reg[59][5]  ( .D(\row2_buffer[60][5] ), .CK(clk), .Q(
        \row2_buffer[59][5] ) );
  DFFQXL \row2_buffer_reg[58][5]  ( .D(\row2_buffer[59][5] ), .CK(clk), .Q(
        \row2_buffer[58][5] ) );
  DFFQXL \row2_buffer_reg[57][5]  ( .D(\row2_buffer[58][5] ), .CK(clk), .Q(
        \row2_buffer[57][5] ) );
  DFFQXL \row2_buffer_reg[56][5]  ( .D(\row2_buffer[57][5] ), .CK(clk), .Q(
        \row2_buffer[56][5] ) );
  DFFQXL \row2_buffer_reg[55][5]  ( .D(\row2_buffer[56][5] ), .CK(clk), .Q(
        \row2_buffer[55][5] ) );
  DFFQXL \row2_buffer_reg[54][5]  ( .D(\row2_buffer[55][5] ), .CK(clk), .Q(
        \row2_buffer[54][5] ) );
  DFFQXL \row2_buffer_reg[53][5]  ( .D(\row2_buffer[54][5] ), .CK(clk), .Q(
        \row2_buffer[53][5] ) );
  DFFQXL \row2_buffer_reg[52][5]  ( .D(\row2_buffer[53][5] ), .CK(clk), .Q(
        \row2_buffer[52][5] ) );
  DFFQXL \row2_buffer_reg[51][5]  ( .D(\row2_buffer[52][5] ), .CK(clk), .Q(
        \row2_buffer[51][5] ) );
  DFFQXL \row2_buffer_reg[50][5]  ( .D(\row2_buffer[51][5] ), .CK(clk), .Q(
        \row2_buffer[50][5] ) );
  DFFQXL \row2_buffer_reg[49][5]  ( .D(\row2_buffer[50][5] ), .CK(clk), .Q(
        \row2_buffer[49][5] ) );
  DFFQXL \row2_buffer_reg[48][5]  ( .D(\row2_buffer[49][5] ), .CK(clk), .Q(
        \row2_buffer[48][5] ) );
  DFFQXL \row2_buffer_reg[47][5]  ( .D(\row2_buffer[48][5] ), .CK(clk), .Q(
        \row2_buffer[47][5] ) );
  DFFQXL \row2_buffer_reg[46][5]  ( .D(\row2_buffer[47][5] ), .CK(clk), .Q(
        \row2_buffer[46][5] ) );
  DFFQXL \row2_buffer_reg[45][5]  ( .D(\row2_buffer[46][5] ), .CK(clk), .Q(
        \row2_buffer[45][5] ) );
  DFFQXL \row2_buffer_reg[44][5]  ( .D(\row2_buffer[45][5] ), .CK(clk), .Q(
        \row2_buffer[44][5] ) );
  DFFQXL \row2_buffer_reg[43][5]  ( .D(\row2_buffer[44][5] ), .CK(clk), .Q(
        \row2_buffer[43][5] ) );
  DFFQXL \row2_buffer_reg[42][5]  ( .D(\row2_buffer[43][5] ), .CK(clk), .Q(
        \row2_buffer[42][5] ) );
  DFFQXL \row2_buffer_reg[41][5]  ( .D(\row2_buffer[42][5] ), .CK(clk), .Q(
        \row2_buffer[41][5] ) );
  DFFQXL \row2_buffer_reg[40][5]  ( .D(\row2_buffer[41][5] ), .CK(clk), .Q(
        \row2_buffer[40][5] ) );
  DFFQXL \row2_buffer_reg[39][5]  ( .D(\row2_buffer[40][5] ), .CK(clk), .Q(
        \row2_buffer[39][5] ) );
  DFFQXL \row2_buffer_reg[38][5]  ( .D(\row2_buffer[39][5] ), .CK(clk), .Q(
        \row2_buffer[38][5] ) );
  DFFQXL \row2_buffer_reg[37][5]  ( .D(\row2_buffer[38][5] ), .CK(clk), .Q(
        \row2_buffer[37][5] ) );
  DFFQXL \row2_buffer_reg[36][5]  ( .D(\row2_buffer[37][5] ), .CK(clk), .Q(
        \row2_buffer[36][5] ) );
  DFFQXL \row2_buffer_reg[35][5]  ( .D(\row2_buffer[36][5] ), .CK(clk), .Q(
        \row2_buffer[35][5] ) );
  DFFQXL \row2_buffer_reg[34][5]  ( .D(\row2_buffer[35][5] ), .CK(clk), .Q(
        \row2_buffer[34][5] ) );
  DFFQXL \row2_buffer_reg[33][5]  ( .D(\row2_buffer[34][5] ), .CK(clk), .Q(
        \row2_buffer[33][5] ) );
  DFFQXL \row2_buffer_reg[32][5]  ( .D(\row2_buffer[33][5] ), .CK(clk), .Q(
        \row2_buffer[32][5] ) );
  DFFQXL \row2_buffer_reg[31][5]  ( .D(\row2_buffer[32][5] ), .CK(clk), .Q(
        \row2_buffer[31][5] ) );
  DFFQXL \row2_buffer_reg[30][5]  ( .D(\row2_buffer[31][5] ), .CK(clk), .Q(
        \row2_buffer[30][5] ) );
  DFFQXL \row2_buffer_reg[29][5]  ( .D(\row2_buffer[30][5] ), .CK(clk), .Q(
        \row2_buffer[29][5] ) );
  DFFQXL \row2_buffer_reg[28][5]  ( .D(\row2_buffer[29][5] ), .CK(clk), .Q(
        \row2_buffer[28][5] ) );
  DFFQXL \row2_buffer_reg[27][5]  ( .D(\row2_buffer[28][5] ), .CK(clk), .Q(
        \row2_buffer[27][5] ) );
  DFFQXL \row2_buffer_reg[26][5]  ( .D(\row2_buffer[27][5] ), .CK(clk), .Q(
        \row2_buffer[26][5] ) );
  DFFQXL \row2_buffer_reg[25][5]  ( .D(\row2_buffer[26][5] ), .CK(clk), .Q(
        \row2_buffer[25][5] ) );
  DFFQXL \row2_buffer_reg[24][5]  ( .D(\row2_buffer[25][5] ), .CK(clk), .Q(
        \row2_buffer[24][5] ) );
  DFFQXL \row2_buffer_reg[23][5]  ( .D(\row2_buffer[24][5] ), .CK(clk), .Q(
        \row2_buffer[23][5] ) );
  DFFQXL \row2_buffer_reg[22][5]  ( .D(\row2_buffer[23][5] ), .CK(clk), .Q(
        \row2_buffer[22][5] ) );
  DFFQXL \row2_buffer_reg[21][5]  ( .D(\row2_buffer[22][5] ), .CK(clk), .Q(
        \row2_buffer[21][5] ) );
  DFFQXL \row2_buffer_reg[20][5]  ( .D(\row2_buffer[21][5] ), .CK(clk), .Q(
        \row2_buffer[20][5] ) );
  DFFQXL \row2_buffer_reg[19][5]  ( .D(\row2_buffer[20][5] ), .CK(clk), .Q(
        \row2_buffer[19][5] ) );
  DFFQXL \row2_buffer_reg[18][5]  ( .D(\row2_buffer[19][5] ), .CK(clk), .Q(
        \row2_buffer[18][5] ) );
  DFFQXL \row2_buffer_reg[17][5]  ( .D(\row2_buffer[18][5] ), .CK(clk), .Q(
        \row2_buffer[17][5] ) );
  DFFQXL \row2_buffer_reg[16][5]  ( .D(\row2_buffer[17][5] ), .CK(clk), .Q(
        \row2_buffer[16][5] ) );
  DFFQXL \row2_buffer_reg[15][5]  ( .D(\row2_buffer[16][5] ), .CK(clk), .Q(
        \row2_buffer[15][5] ) );
  DFFQXL \row2_buffer_reg[14][5]  ( .D(\row2_buffer[15][5] ), .CK(clk), .Q(
        \row2_buffer[14][5] ) );
  DFFQXL \row2_buffer_reg[13][5]  ( .D(\row2_buffer[14][5] ), .CK(clk), .Q(
        \row2_buffer[13][5] ) );
  DFFQXL \row2_buffer_reg[12][5]  ( .D(\row2_buffer[13][5] ), .CK(clk), .Q(
        \row2_buffer[12][5] ) );
  DFFQXL \row2_buffer_reg[11][5]  ( .D(\row2_buffer[12][5] ), .CK(clk), .Q(
        \row2_buffer[11][5] ) );
  DFFQXL \row2_buffer_reg[10][5]  ( .D(\row2_buffer[11][5] ), .CK(clk), .Q(
        \row2_buffer[10][5] ) );
  DFFQXL \row2_buffer_reg[9][5]  ( .D(\row2_buffer[10][5] ), .CK(clk), .Q(
        \row2_buffer[9][5] ) );
  DFFQXL \row2_buffer_reg[8][5]  ( .D(\row2_buffer[9][5] ), .CK(clk), .Q(
        \row2_buffer[8][5] ) );
  DFFQXL \row2_buffer_reg[7][5]  ( .D(\row2_buffer[8][5] ), .CK(clk), .Q(
        \row2_buffer[7][5] ) );
  DFFQXL \row2_buffer_reg[6][5]  ( .D(\row2_buffer[7][5] ), .CK(clk), .Q(
        \row2_buffer[6][5] ) );
  DFFQXL \row2_buffer_reg[5][5]  ( .D(\row2_buffer[6][5] ), .CK(clk), .Q(
        \row2_buffer[5][5] ) );
  DFFQXL \row2_buffer_reg[4][5]  ( .D(\row2_buffer[5][5] ), .CK(clk), .Q(
        \row2_buffer[4][5] ) );
  DFFQXL \row2_buffer_reg[3][5]  ( .D(\row2_buffer[4][5] ), .CK(clk), .Q(
        \row2_buffer[3][5] ) );
  DFFQXL \row1_buffer_reg[225][5]  ( .D(\row2_buffer[0][5] ), .CK(clk), .Q(
        \row1_buffer[225][5] ) );
  DFFQXL \row1_buffer_reg[224][5]  ( .D(\row1_buffer[225][5] ), .CK(clk), .Q(
        \row1_buffer[224][5] ) );
  DFFQXL \row1_buffer_reg[223][5]  ( .D(\row1_buffer[224][5] ), .CK(clk), .Q(
        \row1_buffer[223][5] ) );
  DFFQXL \row1_buffer_reg[222][5]  ( .D(\row1_buffer[223][5] ), .CK(clk), .Q(
        \row1_buffer[222][5] ) );
  DFFQXL \row1_buffer_reg[221][5]  ( .D(\row1_buffer[222][5] ), .CK(clk), .Q(
        \row1_buffer[221][5] ) );
  DFFQXL \row1_buffer_reg[220][5]  ( .D(\row1_buffer[221][5] ), .CK(clk), .Q(
        \row1_buffer[220][5] ) );
  DFFQXL \row1_buffer_reg[219][5]  ( .D(\row1_buffer[220][5] ), .CK(clk), .Q(
        \row1_buffer[219][5] ) );
  DFFQXL \row1_buffer_reg[218][5]  ( .D(\row1_buffer[219][5] ), .CK(clk), .Q(
        \row1_buffer[218][5] ) );
  DFFQXL \row1_buffer_reg[217][5]  ( .D(\row1_buffer[218][5] ), .CK(clk), .Q(
        \row1_buffer[217][5] ) );
  DFFQXL \row1_buffer_reg[216][5]  ( .D(\row1_buffer[217][5] ), .CK(clk), .Q(
        \row1_buffer[216][5] ) );
  DFFQXL \row1_buffer_reg[215][5]  ( .D(\row1_buffer[216][5] ), .CK(clk), .Q(
        \row1_buffer[215][5] ) );
  DFFQXL \row1_buffer_reg[214][5]  ( .D(\row1_buffer[215][5] ), .CK(clk), .Q(
        \row1_buffer[214][5] ) );
  DFFQXL \row1_buffer_reg[213][5]  ( .D(\row1_buffer[214][5] ), .CK(clk), .Q(
        \row1_buffer[213][5] ) );
  DFFQXL \row1_buffer_reg[212][5]  ( .D(\row1_buffer[213][5] ), .CK(clk), .Q(
        \row1_buffer[212][5] ) );
  DFFQXL \row1_buffer_reg[211][5]  ( .D(\row1_buffer[212][5] ), .CK(clk), .Q(
        \row1_buffer[211][5] ) );
  DFFQXL \row1_buffer_reg[210][5]  ( .D(\row1_buffer[211][5] ), .CK(clk), .Q(
        \row1_buffer[210][5] ) );
  DFFQXL \row1_buffer_reg[209][5]  ( .D(\row1_buffer[210][5] ), .CK(clk), .Q(
        \row1_buffer[209][5] ) );
  DFFQXL \row1_buffer_reg[208][5]  ( .D(\row1_buffer[209][5] ), .CK(clk), .Q(
        \row1_buffer[208][5] ) );
  DFFQXL \row1_buffer_reg[207][5]  ( .D(\row1_buffer[208][5] ), .CK(clk), .Q(
        \row1_buffer[207][5] ) );
  DFFQXL \row1_buffer_reg[206][5]  ( .D(\row1_buffer[207][5] ), .CK(clk), .Q(
        \row1_buffer[206][5] ) );
  DFFQXL \row1_buffer_reg[205][5]  ( .D(\row1_buffer[206][5] ), .CK(clk), .Q(
        \row1_buffer[205][5] ) );
  DFFQXL \row1_buffer_reg[204][5]  ( .D(\row1_buffer[205][5] ), .CK(clk), .Q(
        \row1_buffer[204][5] ) );
  DFFQXL \row1_buffer_reg[203][5]  ( .D(\row1_buffer[204][5] ), .CK(clk), .Q(
        \row1_buffer[203][5] ) );
  DFFQXL \row1_buffer_reg[202][5]  ( .D(\row1_buffer[203][5] ), .CK(clk), .Q(
        \row1_buffer[202][5] ) );
  DFFQXL \row1_buffer_reg[201][5]  ( .D(\row1_buffer[202][5] ), .CK(clk), .Q(
        \row1_buffer[201][5] ) );
  DFFQXL \row1_buffer_reg[200][5]  ( .D(\row1_buffer[201][5] ), .CK(clk), .Q(
        \row1_buffer[200][5] ) );
  DFFQXL \row1_buffer_reg[199][5]  ( .D(\row1_buffer[200][5] ), .CK(clk), .Q(
        \row1_buffer[199][5] ) );
  DFFQXL \row1_buffer_reg[198][5]  ( .D(\row1_buffer[199][5] ), .CK(clk), .Q(
        \row1_buffer[198][5] ) );
  DFFQXL \row1_buffer_reg[197][5]  ( .D(\row1_buffer[198][5] ), .CK(clk), .Q(
        \row1_buffer[197][5] ) );
  DFFQXL \row1_buffer_reg[196][5]  ( .D(\row1_buffer[197][5] ), .CK(clk), .Q(
        \row1_buffer[196][5] ) );
  DFFQXL \row1_buffer_reg[195][5]  ( .D(\row1_buffer[196][5] ), .CK(clk), .Q(
        \row1_buffer[195][5] ) );
  DFFQXL \row1_buffer_reg[194][5]  ( .D(\row1_buffer[195][5] ), .CK(clk), .Q(
        \row1_buffer[194][5] ) );
  DFFQXL \row1_buffer_reg[193][5]  ( .D(\row1_buffer[194][5] ), .CK(clk), .Q(
        \row1_buffer[193][5] ) );
  DFFQXL \row1_buffer_reg[192][5]  ( .D(\row1_buffer[193][5] ), .CK(clk), .Q(
        \row1_buffer[192][5] ) );
  DFFQXL \row1_buffer_reg[191][5]  ( .D(\row1_buffer[192][5] ), .CK(clk), .Q(
        \row1_buffer[191][5] ) );
  DFFQXL \row1_buffer_reg[190][5]  ( .D(\row1_buffer[191][5] ), .CK(clk), .Q(
        \row1_buffer[190][5] ) );
  DFFQXL \row1_buffer_reg[189][5]  ( .D(\row1_buffer[190][5] ), .CK(clk), .Q(
        \row1_buffer[189][5] ) );
  DFFQXL \row1_buffer_reg[188][5]  ( .D(\row1_buffer[189][5] ), .CK(clk), .Q(
        \row1_buffer[188][5] ) );
  DFFQXL \row1_buffer_reg[187][5]  ( .D(\row1_buffer[188][5] ), .CK(clk), .Q(
        \row1_buffer[187][5] ) );
  DFFQXL \row1_buffer_reg[186][5]  ( .D(\row1_buffer[187][5] ), .CK(clk), .Q(
        \row1_buffer[186][5] ) );
  DFFQXL \row1_buffer_reg[185][5]  ( .D(\row1_buffer[186][5] ), .CK(clk), .Q(
        \row1_buffer[185][5] ) );
  DFFQXL \row1_buffer_reg[184][5]  ( .D(\row1_buffer[185][5] ), .CK(clk), .Q(
        \row1_buffer[184][5] ) );
  DFFQXL \row1_buffer_reg[183][5]  ( .D(\row1_buffer[184][5] ), .CK(clk), .Q(
        \row1_buffer[183][5] ) );
  DFFQXL \row1_buffer_reg[182][5]  ( .D(\row1_buffer[183][5] ), .CK(clk), .Q(
        \row1_buffer[182][5] ) );
  DFFQXL \row1_buffer_reg[181][5]  ( .D(\row1_buffer[182][5] ), .CK(clk), .Q(
        \row1_buffer[181][5] ) );
  DFFQXL \row1_buffer_reg[180][5]  ( .D(\row1_buffer[181][5] ), .CK(clk), .Q(
        \row1_buffer[180][5] ) );
  DFFQXL \row1_buffer_reg[179][5]  ( .D(\row1_buffer[180][5] ), .CK(clk), .Q(
        \row1_buffer[179][5] ) );
  DFFQXL \row1_buffer_reg[178][5]  ( .D(\row1_buffer[179][5] ), .CK(clk), .Q(
        \row1_buffer[178][5] ) );
  DFFQXL \row1_buffer_reg[177][5]  ( .D(\row1_buffer[178][5] ), .CK(clk), .Q(
        \row1_buffer[177][5] ) );
  DFFQXL \row1_buffer_reg[176][5]  ( .D(\row1_buffer[177][5] ), .CK(clk), .Q(
        \row1_buffer[176][5] ) );
  DFFQXL \row1_buffer_reg[175][5]  ( .D(\row1_buffer[176][5] ), .CK(clk), .Q(
        \row1_buffer[175][5] ) );
  DFFQXL \row1_buffer_reg[174][5]  ( .D(\row1_buffer[175][5] ), .CK(clk), .Q(
        \row1_buffer[174][5] ) );
  DFFQXL \row1_buffer_reg[173][5]  ( .D(\row1_buffer[174][5] ), .CK(clk), .Q(
        \row1_buffer[173][5] ) );
  DFFQXL \row1_buffer_reg[172][5]  ( .D(\row1_buffer[173][5] ), .CK(clk), .Q(
        \row1_buffer[172][5] ) );
  DFFQXL \row1_buffer_reg[171][5]  ( .D(\row1_buffer[172][5] ), .CK(clk), .Q(
        \row1_buffer[171][5] ) );
  DFFQXL \row1_buffer_reg[170][5]  ( .D(\row1_buffer[171][5] ), .CK(clk), .Q(
        \row1_buffer[170][5] ) );
  DFFQXL \row1_buffer_reg[169][5]  ( .D(\row1_buffer[170][5] ), .CK(clk), .Q(
        \row1_buffer[169][5] ) );
  DFFQXL \row1_buffer_reg[168][5]  ( .D(\row1_buffer[169][5] ), .CK(clk), .Q(
        \row1_buffer[168][5] ) );
  DFFQXL \row1_buffer_reg[167][5]  ( .D(\row1_buffer[168][5] ), .CK(clk), .Q(
        \row1_buffer[167][5] ) );
  DFFQXL \row1_buffer_reg[166][5]  ( .D(\row1_buffer[167][5] ), .CK(clk), .Q(
        \row1_buffer[166][5] ) );
  DFFQXL \row1_buffer_reg[165][5]  ( .D(\row1_buffer[166][5] ), .CK(clk), .Q(
        \row1_buffer[165][5] ) );
  DFFQXL \row1_buffer_reg[164][5]  ( .D(\row1_buffer[165][5] ), .CK(clk), .Q(
        \row1_buffer[164][5] ) );
  DFFQXL \row1_buffer_reg[163][5]  ( .D(\row1_buffer[164][5] ), .CK(clk), .Q(
        \row1_buffer[163][5] ) );
  DFFQXL \row1_buffer_reg[162][5]  ( .D(\row1_buffer[163][5] ), .CK(clk), .Q(
        \row1_buffer[162][5] ) );
  DFFQXL \row1_buffer_reg[161][5]  ( .D(\row1_buffer[162][5] ), .CK(clk), .Q(
        \row1_buffer[161][5] ) );
  DFFQXL \row1_buffer_reg[160][5]  ( .D(\row1_buffer[161][5] ), .CK(clk), .Q(
        \row1_buffer[160][5] ) );
  DFFQXL \row1_buffer_reg[159][5]  ( .D(\row1_buffer[160][5] ), .CK(clk), .Q(
        \row1_buffer[159][5] ) );
  DFFQXL \row1_buffer_reg[158][5]  ( .D(\row1_buffer[159][5] ), .CK(clk), .Q(
        \row1_buffer[158][5] ) );
  DFFQXL \row1_buffer_reg[157][5]  ( .D(\row1_buffer[158][5] ), .CK(clk), .Q(
        \row1_buffer[157][5] ) );
  DFFQXL \row1_buffer_reg[156][5]  ( .D(\row1_buffer[157][5] ), .CK(clk), .Q(
        \row1_buffer[156][5] ) );
  DFFQXL \row1_buffer_reg[155][5]  ( .D(\row1_buffer[156][5] ), .CK(clk), .Q(
        \row1_buffer[155][5] ) );
  DFFQXL \row1_buffer_reg[154][5]  ( .D(\row1_buffer[155][5] ), .CK(clk), .Q(
        \row1_buffer[154][5] ) );
  DFFQXL \row1_buffer_reg[153][5]  ( .D(\row1_buffer[154][5] ), .CK(clk), .Q(
        \row1_buffer[153][5] ) );
  DFFQXL \row1_buffer_reg[152][5]  ( .D(\row1_buffer[153][5] ), .CK(clk), .Q(
        \row1_buffer[152][5] ) );
  DFFQXL \row1_buffer_reg[151][5]  ( .D(\row1_buffer[152][5] ), .CK(clk), .Q(
        \row1_buffer[151][5] ) );
  DFFQXL \row1_buffer_reg[150][5]  ( .D(\row1_buffer[151][5] ), .CK(clk), .Q(
        \row1_buffer[150][5] ) );
  DFFQXL \row1_buffer_reg[149][5]  ( .D(\row1_buffer[150][5] ), .CK(clk), .Q(
        \row1_buffer[149][5] ) );
  DFFQXL \row1_buffer_reg[148][5]  ( .D(\row1_buffer[149][5] ), .CK(clk), .Q(
        \row1_buffer[148][5] ) );
  DFFQXL \row1_buffer_reg[147][5]  ( .D(\row1_buffer[148][5] ), .CK(clk), .Q(
        \row1_buffer[147][5] ) );
  DFFQXL \row1_buffer_reg[146][5]  ( .D(\row1_buffer[147][5] ), .CK(clk), .Q(
        \row1_buffer[146][5] ) );
  DFFQXL \row1_buffer_reg[145][5]  ( .D(\row1_buffer[146][5] ), .CK(clk), .Q(
        \row1_buffer[145][5] ) );
  DFFQXL \row1_buffer_reg[144][5]  ( .D(\row1_buffer[145][5] ), .CK(clk), .Q(
        \row1_buffer[144][5] ) );
  DFFQXL \row1_buffer_reg[143][5]  ( .D(\row1_buffer[144][5] ), .CK(clk), .Q(
        \row1_buffer[143][5] ) );
  DFFQXL \row1_buffer_reg[142][5]  ( .D(\row1_buffer[143][5] ), .CK(clk), .Q(
        \row1_buffer[142][5] ) );
  DFFQXL \row1_buffer_reg[141][5]  ( .D(\row1_buffer[142][5] ), .CK(clk), .Q(
        \row1_buffer[141][5] ) );
  DFFQXL \row1_buffer_reg[140][5]  ( .D(\row1_buffer[141][5] ), .CK(clk), .Q(
        \row1_buffer[140][5] ) );
  DFFQXL \row1_buffer_reg[139][5]  ( .D(\row1_buffer[140][5] ), .CK(clk), .Q(
        \row1_buffer[139][5] ) );
  DFFQXL \row1_buffer_reg[138][5]  ( .D(\row1_buffer[139][5] ), .CK(clk), .Q(
        \row1_buffer[138][5] ) );
  DFFQXL \row1_buffer_reg[137][5]  ( .D(\row1_buffer[138][5] ), .CK(clk), .Q(
        \row1_buffer[137][5] ) );
  DFFQXL \row1_buffer_reg[136][5]  ( .D(\row1_buffer[137][5] ), .CK(clk), .Q(
        \row1_buffer[136][5] ) );
  DFFQXL \row1_buffer_reg[135][5]  ( .D(\row1_buffer[136][5] ), .CK(clk), .Q(
        \row1_buffer[135][5] ) );
  DFFQXL \row1_buffer_reg[134][5]  ( .D(\row1_buffer[135][5] ), .CK(clk), .Q(
        \row1_buffer[134][5] ) );
  DFFQXL \row1_buffer_reg[133][5]  ( .D(\row1_buffer[134][5] ), .CK(clk), .Q(
        \row1_buffer[133][5] ) );
  DFFQXL \row1_buffer_reg[132][5]  ( .D(\row1_buffer[133][5] ), .CK(clk), .Q(
        \row1_buffer[132][5] ) );
  DFFQXL \row1_buffer_reg[131][5]  ( .D(\row1_buffer[132][5] ), .CK(clk), .Q(
        \row1_buffer[131][5] ) );
  DFFQXL \row1_buffer_reg[130][5]  ( .D(\row1_buffer[131][5] ), .CK(clk), .Q(
        \row1_buffer[130][5] ) );
  DFFQXL \row1_buffer_reg[129][5]  ( .D(\row1_buffer[130][5] ), .CK(clk), .Q(
        \row1_buffer[129][5] ) );
  DFFQXL \row1_buffer_reg[128][5]  ( .D(\row1_buffer[129][5] ), .CK(clk), .Q(
        \row1_buffer[128][5] ) );
  DFFQXL \row1_buffer_reg[127][5]  ( .D(\row1_buffer[128][5] ), .CK(clk), .Q(
        \row1_buffer[127][5] ) );
  DFFQXL \row1_buffer_reg[126][5]  ( .D(\row1_buffer[127][5] ), .CK(clk), .Q(
        \row1_buffer[126][5] ) );
  DFFQXL \row1_buffer_reg[125][5]  ( .D(\row1_buffer[126][5] ), .CK(clk), .Q(
        \row1_buffer[125][5] ) );
  DFFQXL \row1_buffer_reg[124][5]  ( .D(\row1_buffer[125][5] ), .CK(clk), .Q(
        \row1_buffer[124][5] ) );
  DFFQXL \row1_buffer_reg[123][5]  ( .D(\row1_buffer[124][5] ), .CK(clk), .Q(
        \row1_buffer[123][5] ) );
  DFFQXL \row1_buffer_reg[122][5]  ( .D(\row1_buffer[123][5] ), .CK(clk), .Q(
        \row1_buffer[122][5] ) );
  DFFQXL \row1_buffer_reg[121][5]  ( .D(\row1_buffer[122][5] ), .CK(clk), .Q(
        \row1_buffer[121][5] ) );
  DFFQXL \row1_buffer_reg[120][5]  ( .D(\row1_buffer[121][5] ), .CK(clk), .Q(
        \row1_buffer[120][5] ) );
  DFFQXL \row1_buffer_reg[119][5]  ( .D(\row1_buffer[120][5] ), .CK(clk), .Q(
        \row1_buffer[119][5] ) );
  DFFQXL \row1_buffer_reg[118][5]  ( .D(\row1_buffer[119][5] ), .CK(clk), .Q(
        \row1_buffer[118][5] ) );
  DFFQXL \row1_buffer_reg[117][5]  ( .D(\row1_buffer[118][5] ), .CK(clk), .Q(
        \row1_buffer[117][5] ) );
  DFFQXL \row1_buffer_reg[116][5]  ( .D(\row1_buffer[117][5] ), .CK(clk), .Q(
        \row1_buffer[116][5] ) );
  DFFQXL \row1_buffer_reg[115][5]  ( .D(\row1_buffer[116][5] ), .CK(clk), .Q(
        \row1_buffer[115][5] ) );
  DFFQXL \row1_buffer_reg[114][5]  ( .D(\row1_buffer[115][5] ), .CK(clk), .Q(
        \row1_buffer[114][5] ) );
  DFFQXL \row1_buffer_reg[113][5]  ( .D(\row1_buffer[114][5] ), .CK(clk), .Q(
        \row1_buffer[113][5] ) );
  DFFQXL \row1_buffer_reg[112][5]  ( .D(\row1_buffer[113][5] ), .CK(clk), .Q(
        \row1_buffer[112][5] ) );
  DFFQXL \row1_buffer_reg[111][5]  ( .D(\row1_buffer[112][5] ), .CK(clk), .Q(
        \row1_buffer[111][5] ) );
  DFFQXL \row1_buffer_reg[110][5]  ( .D(\row1_buffer[111][5] ), .CK(clk), .Q(
        \row1_buffer[110][5] ) );
  DFFQXL \row1_buffer_reg[109][5]  ( .D(\row1_buffer[110][5] ), .CK(clk), .Q(
        \row1_buffer[109][5] ) );
  DFFQXL \row1_buffer_reg[108][5]  ( .D(\row1_buffer[109][5] ), .CK(clk), .Q(
        \row1_buffer[108][5] ) );
  DFFQXL \row1_buffer_reg[107][5]  ( .D(\row1_buffer[108][5] ), .CK(clk), .Q(
        \row1_buffer[107][5] ) );
  DFFQXL \row1_buffer_reg[106][5]  ( .D(\row1_buffer[107][5] ), .CK(clk), .Q(
        \row1_buffer[106][5] ) );
  DFFQXL \row1_buffer_reg[105][5]  ( .D(\row1_buffer[106][5] ), .CK(clk), .Q(
        \row1_buffer[105][5] ) );
  DFFQXL \row1_buffer_reg[104][5]  ( .D(\row1_buffer[105][5] ), .CK(clk), .Q(
        \row1_buffer[104][5] ) );
  DFFQXL \row1_buffer_reg[103][5]  ( .D(\row1_buffer[104][5] ), .CK(clk), .Q(
        \row1_buffer[103][5] ) );
  DFFQXL \row1_buffer_reg[102][5]  ( .D(\row1_buffer[103][5] ), .CK(clk), .Q(
        \row1_buffer[102][5] ) );
  DFFQXL \row1_buffer_reg[101][5]  ( .D(\row1_buffer[102][5] ), .CK(clk), .Q(
        \row1_buffer[101][5] ) );
  DFFQXL \row1_buffer_reg[100][5]  ( .D(\row1_buffer[101][5] ), .CK(clk), .Q(
        \row1_buffer[100][5] ) );
  DFFQXL \row1_buffer_reg[99][5]  ( .D(\row1_buffer[100][5] ), .CK(clk), .Q(
        \row1_buffer[99][5] ) );
  DFFQXL \row1_buffer_reg[98][5]  ( .D(\row1_buffer[99][5] ), .CK(clk), .Q(
        \row1_buffer[98][5] ) );
  DFFQXL \row1_buffer_reg[97][5]  ( .D(\row1_buffer[98][5] ), .CK(clk), .Q(
        \row1_buffer[97][5] ) );
  DFFQXL \row1_buffer_reg[96][5]  ( .D(\row1_buffer[97][5] ), .CK(clk), .Q(
        \row1_buffer[96][5] ) );
  DFFQXL \row1_buffer_reg[95][5]  ( .D(\row1_buffer[96][5] ), .CK(clk), .Q(
        \row1_buffer[95][5] ) );
  DFFQXL \row1_buffer_reg[94][5]  ( .D(\row1_buffer[95][5] ), .CK(clk), .Q(
        \row1_buffer[94][5] ) );
  DFFQXL \row1_buffer_reg[93][5]  ( .D(\row1_buffer[94][5] ), .CK(clk), .Q(
        \row1_buffer[93][5] ) );
  DFFQXL \row1_buffer_reg[92][5]  ( .D(\row1_buffer[93][5] ), .CK(clk), .Q(
        \row1_buffer[92][5] ) );
  DFFQXL \row1_buffer_reg[91][5]  ( .D(\row1_buffer[92][5] ), .CK(clk), .Q(
        \row1_buffer[91][5] ) );
  DFFQXL \row1_buffer_reg[90][5]  ( .D(\row1_buffer[91][5] ), .CK(clk), .Q(
        \row1_buffer[90][5] ) );
  DFFQXL \row1_buffer_reg[89][5]  ( .D(\row1_buffer[90][5] ), .CK(clk), .Q(
        \row1_buffer[89][5] ) );
  DFFQXL \row1_buffer_reg[88][5]  ( .D(\row1_buffer[89][5] ), .CK(clk), .Q(
        \row1_buffer[88][5] ) );
  DFFQXL \row1_buffer_reg[87][5]  ( .D(\row1_buffer[88][5] ), .CK(clk), .Q(
        \row1_buffer[87][5] ) );
  DFFQXL \row1_buffer_reg[86][5]  ( .D(\row1_buffer[87][5] ), .CK(clk), .Q(
        \row1_buffer[86][5] ) );
  DFFQXL \row1_buffer_reg[85][5]  ( .D(\row1_buffer[86][5] ), .CK(clk), .Q(
        \row1_buffer[85][5] ) );
  DFFQXL \row1_buffer_reg[84][5]  ( .D(\row1_buffer[85][5] ), .CK(clk), .Q(
        \row1_buffer[84][5] ) );
  DFFQXL \row1_buffer_reg[83][5]  ( .D(\row1_buffer[84][5] ), .CK(clk), .Q(
        \row1_buffer[83][5] ) );
  DFFQXL \row1_buffer_reg[82][5]  ( .D(\row1_buffer[83][5] ), .CK(clk), .Q(
        \row1_buffer[82][5] ) );
  DFFQXL \row1_buffer_reg[81][5]  ( .D(\row1_buffer[82][5] ), .CK(clk), .Q(
        \row1_buffer[81][5] ) );
  DFFQXL \row1_buffer_reg[80][5]  ( .D(\row1_buffer[81][5] ), .CK(clk), .Q(
        \row1_buffer[80][5] ) );
  DFFQXL \row1_buffer_reg[79][5]  ( .D(\row1_buffer[80][5] ), .CK(clk), .Q(
        \row1_buffer[79][5] ) );
  DFFQXL \row1_buffer_reg[78][5]  ( .D(\row1_buffer[79][5] ), .CK(clk), .Q(
        \row1_buffer[78][5] ) );
  DFFQXL \row1_buffer_reg[77][5]  ( .D(\row1_buffer[78][5] ), .CK(clk), .Q(
        \row1_buffer[77][5] ) );
  DFFQXL \row1_buffer_reg[76][5]  ( .D(\row1_buffer[77][5] ), .CK(clk), .Q(
        \row1_buffer[76][5] ) );
  DFFQXL \row1_buffer_reg[75][5]  ( .D(\row1_buffer[76][5] ), .CK(clk), .Q(
        \row1_buffer[75][5] ) );
  DFFQXL \row1_buffer_reg[74][5]  ( .D(\row1_buffer[75][5] ), .CK(clk), .Q(
        \row1_buffer[74][5] ) );
  DFFQXL \row1_buffer_reg[73][5]  ( .D(\row1_buffer[74][5] ), .CK(clk), .Q(
        \row1_buffer[73][5] ) );
  DFFQXL \row1_buffer_reg[72][5]  ( .D(\row1_buffer[73][5] ), .CK(clk), .Q(
        \row1_buffer[72][5] ) );
  DFFQXL \row1_buffer_reg[71][5]  ( .D(\row1_buffer[72][5] ), .CK(clk), .Q(
        \row1_buffer[71][5] ) );
  DFFQXL \row1_buffer_reg[70][5]  ( .D(\row1_buffer[71][5] ), .CK(clk), .Q(
        \row1_buffer[70][5] ) );
  DFFQXL \row1_buffer_reg[69][5]  ( .D(\row1_buffer[70][5] ), .CK(clk), .Q(
        \row1_buffer[69][5] ) );
  DFFQXL \row1_buffer_reg[68][5]  ( .D(\row1_buffer[69][5] ), .CK(clk), .Q(
        \row1_buffer[68][5] ) );
  DFFQXL \row1_buffer_reg[67][5]  ( .D(\row1_buffer[68][5] ), .CK(clk), .Q(
        \row1_buffer[67][5] ) );
  DFFQXL \row1_buffer_reg[66][5]  ( .D(\row1_buffer[67][5] ), .CK(clk), .Q(
        \row1_buffer[66][5] ) );
  DFFQXL \row1_buffer_reg[65][5]  ( .D(\row1_buffer[66][5] ), .CK(clk), .Q(
        \row1_buffer[65][5] ) );
  DFFQXL \row1_buffer_reg[64][5]  ( .D(\row1_buffer[65][5] ), .CK(clk), .Q(
        \row1_buffer[64][5] ) );
  DFFQXL \row1_buffer_reg[63][5]  ( .D(\row1_buffer[64][5] ), .CK(clk), .Q(
        \row1_buffer[63][5] ) );
  DFFQXL \row1_buffer_reg[62][5]  ( .D(\row1_buffer[63][5] ), .CK(clk), .Q(
        \row1_buffer[62][5] ) );
  DFFQXL \row1_buffer_reg[61][5]  ( .D(\row1_buffer[62][5] ), .CK(clk), .Q(
        \row1_buffer[61][5] ) );
  DFFQXL \row1_buffer_reg[60][5]  ( .D(\row1_buffer[61][5] ), .CK(clk), .Q(
        \row1_buffer[60][5] ) );
  DFFQXL \row1_buffer_reg[59][5]  ( .D(\row1_buffer[60][5] ), .CK(clk), .Q(
        \row1_buffer[59][5] ) );
  DFFQXL \row1_buffer_reg[58][5]  ( .D(\row1_buffer[59][5] ), .CK(clk), .Q(
        \row1_buffer[58][5] ) );
  DFFQXL \row1_buffer_reg[57][5]  ( .D(\row1_buffer[58][5] ), .CK(clk), .Q(
        \row1_buffer[57][5] ) );
  DFFQXL \row1_buffer_reg[56][5]  ( .D(\row1_buffer[57][5] ), .CK(clk), .Q(
        \row1_buffer[56][5] ) );
  DFFQXL \row1_buffer_reg[55][5]  ( .D(\row1_buffer[56][5] ), .CK(clk), .Q(
        \row1_buffer[55][5] ) );
  DFFQXL \row1_buffer_reg[54][5]  ( .D(\row1_buffer[55][5] ), .CK(clk), .Q(
        \row1_buffer[54][5] ) );
  DFFQXL \row1_buffer_reg[53][5]  ( .D(\row1_buffer[54][5] ), .CK(clk), .Q(
        \row1_buffer[53][5] ) );
  DFFQXL \row1_buffer_reg[52][5]  ( .D(\row1_buffer[53][5] ), .CK(clk), .Q(
        \row1_buffer[52][5] ) );
  DFFQXL \row1_buffer_reg[51][5]  ( .D(\row1_buffer[52][5] ), .CK(clk), .Q(
        \row1_buffer[51][5] ) );
  DFFQXL \row1_buffer_reg[50][5]  ( .D(\row1_buffer[51][5] ), .CK(clk), .Q(
        \row1_buffer[50][5] ) );
  DFFQXL \row1_buffer_reg[49][5]  ( .D(\row1_buffer[50][5] ), .CK(clk), .Q(
        \row1_buffer[49][5] ) );
  DFFQXL \row1_buffer_reg[48][5]  ( .D(\row1_buffer[49][5] ), .CK(clk), .Q(
        \row1_buffer[48][5] ) );
  DFFQXL \row1_buffer_reg[47][5]  ( .D(\row1_buffer[48][5] ), .CK(clk), .Q(
        \row1_buffer[47][5] ) );
  DFFQXL \row1_buffer_reg[46][5]  ( .D(\row1_buffer[47][5] ), .CK(clk), .Q(
        \row1_buffer[46][5] ) );
  DFFQXL \row1_buffer_reg[45][5]  ( .D(\row1_buffer[46][5] ), .CK(clk), .Q(
        \row1_buffer[45][5] ) );
  DFFQXL \row1_buffer_reg[44][5]  ( .D(\row1_buffer[45][5] ), .CK(clk), .Q(
        \row1_buffer[44][5] ) );
  DFFQXL \row1_buffer_reg[43][5]  ( .D(\row1_buffer[44][5] ), .CK(clk), .Q(
        \row1_buffer[43][5] ) );
  DFFQXL \row1_buffer_reg[42][5]  ( .D(\row1_buffer[43][5] ), .CK(clk), .Q(
        \row1_buffer[42][5] ) );
  DFFQXL \row1_buffer_reg[41][5]  ( .D(\row1_buffer[42][5] ), .CK(clk), .Q(
        \row1_buffer[41][5] ) );
  DFFQXL \row1_buffer_reg[40][5]  ( .D(\row1_buffer[41][5] ), .CK(clk), .Q(
        \row1_buffer[40][5] ) );
  DFFQXL \row1_buffer_reg[39][5]  ( .D(\row1_buffer[40][5] ), .CK(clk), .Q(
        \row1_buffer[39][5] ) );
  DFFQXL \row1_buffer_reg[38][5]  ( .D(\row1_buffer[39][5] ), .CK(clk), .Q(
        \row1_buffer[38][5] ) );
  DFFQXL \row1_buffer_reg[37][5]  ( .D(\row1_buffer[38][5] ), .CK(clk), .Q(
        \row1_buffer[37][5] ) );
  DFFQXL \row1_buffer_reg[36][5]  ( .D(\row1_buffer[37][5] ), .CK(clk), .Q(
        \row1_buffer[36][5] ) );
  DFFQXL \row1_buffer_reg[35][5]  ( .D(\row1_buffer[36][5] ), .CK(clk), .Q(
        \row1_buffer[35][5] ) );
  DFFQXL \row1_buffer_reg[34][5]  ( .D(\row1_buffer[35][5] ), .CK(clk), .Q(
        \row1_buffer[34][5] ) );
  DFFQXL \row1_buffer_reg[33][5]  ( .D(\row1_buffer[34][5] ), .CK(clk), .Q(
        \row1_buffer[33][5] ) );
  DFFQXL \row1_buffer_reg[32][5]  ( .D(\row1_buffer[33][5] ), .CK(clk), .Q(
        \row1_buffer[32][5] ) );
  DFFQXL \row1_buffer_reg[31][5]  ( .D(\row1_buffer[32][5] ), .CK(clk), .Q(
        \row1_buffer[31][5] ) );
  DFFQXL \row1_buffer_reg[30][5]  ( .D(\row1_buffer[31][5] ), .CK(clk), .Q(
        \row1_buffer[30][5] ) );
  DFFQXL \row1_buffer_reg[29][5]  ( .D(\row1_buffer[30][5] ), .CK(clk), .Q(
        \row1_buffer[29][5] ) );
  DFFQXL \row1_buffer_reg[28][5]  ( .D(\row1_buffer[29][5] ), .CK(clk), .Q(
        \row1_buffer[28][5] ) );
  DFFQXL \row1_buffer_reg[27][5]  ( .D(\row1_buffer[28][5] ), .CK(clk), .Q(
        \row1_buffer[27][5] ) );
  DFFQXL \row1_buffer_reg[26][5]  ( .D(\row1_buffer[27][5] ), .CK(clk), .Q(
        \row1_buffer[26][5] ) );
  DFFQXL \row1_buffer_reg[25][5]  ( .D(\row1_buffer[26][5] ), .CK(clk), .Q(
        \row1_buffer[25][5] ) );
  DFFQXL \row1_buffer_reg[24][5]  ( .D(\row1_buffer[25][5] ), .CK(clk), .Q(
        \row1_buffer[24][5] ) );
  DFFQXL \row1_buffer_reg[23][5]  ( .D(\row1_buffer[24][5] ), .CK(clk), .Q(
        \row1_buffer[23][5] ) );
  DFFQXL \row1_buffer_reg[22][5]  ( .D(\row1_buffer[23][5] ), .CK(clk), .Q(
        \row1_buffer[22][5] ) );
  DFFQXL \row1_buffer_reg[21][5]  ( .D(\row1_buffer[22][5] ), .CK(clk), .Q(
        \row1_buffer[21][5] ) );
  DFFQXL \row1_buffer_reg[20][5]  ( .D(\row1_buffer[21][5] ), .CK(clk), .Q(
        \row1_buffer[20][5] ) );
  DFFQXL \row1_buffer_reg[19][5]  ( .D(\row1_buffer[20][5] ), .CK(clk), .Q(
        \row1_buffer[19][5] ) );
  DFFQXL \row1_buffer_reg[18][5]  ( .D(\row1_buffer[19][5] ), .CK(clk), .Q(
        \row1_buffer[18][5] ) );
  DFFQXL \row1_buffer_reg[17][5]  ( .D(\row1_buffer[18][5] ), .CK(clk), .Q(
        \row1_buffer[17][5] ) );
  DFFQXL \row1_buffer_reg[16][5]  ( .D(\row1_buffer[17][5] ), .CK(clk), .Q(
        \row1_buffer[16][5] ) );
  DFFQXL \row1_buffer_reg[15][5]  ( .D(\row1_buffer[16][5] ), .CK(clk), .Q(
        \row1_buffer[15][5] ) );
  DFFQXL \row1_buffer_reg[14][5]  ( .D(\row1_buffer[15][5] ), .CK(clk), .Q(
        \row1_buffer[14][5] ) );
  DFFQXL \row1_buffer_reg[13][5]  ( .D(\row1_buffer[14][5] ), .CK(clk), .Q(
        \row1_buffer[13][5] ) );
  DFFQXL \row1_buffer_reg[12][5]  ( .D(\row1_buffer[13][5] ), .CK(clk), .Q(
        \row1_buffer[12][5] ) );
  DFFQXL \row1_buffer_reg[11][5]  ( .D(\row1_buffer[12][5] ), .CK(clk), .Q(
        \row1_buffer[11][5] ) );
  DFFQXL \row1_buffer_reg[10][5]  ( .D(\row1_buffer[11][5] ), .CK(clk), .Q(
        \row1_buffer[10][5] ) );
  DFFQXL \row1_buffer_reg[9][5]  ( .D(\row1_buffer[10][5] ), .CK(clk), .Q(
        \row1_buffer[9][5] ) );
  DFFQXL \row1_buffer_reg[8][5]  ( .D(\row1_buffer[9][5] ), .CK(clk), .Q(
        \row1_buffer[8][5] ) );
  DFFQXL \row1_buffer_reg[7][5]  ( .D(\row1_buffer[8][5] ), .CK(clk), .Q(
        \row1_buffer[7][5] ) );
  DFFQXL \row1_buffer_reg[6][5]  ( .D(\row1_buffer[7][5] ), .CK(clk), .Q(
        \row1_buffer[6][5] ) );
  DFFQXL \row1_buffer_reg[5][5]  ( .D(\row1_buffer[6][5] ), .CK(clk), .Q(
        \row1_buffer[5][5] ) );
  DFFQXL \row1_buffer_reg[4][5]  ( .D(\row1_buffer[5][5] ), .CK(clk), .Q(
        \row1_buffer[4][5] ) );
  DFFQXL \row1_buffer_reg[3][5]  ( .D(\row1_buffer[4][5] ), .CK(clk), .Q(
        \row1_buffer[3][5] ) );
  DFFQXL \row1_buffer_reg[0][5]  ( .D(\row1_buffer[1][5] ), .CK(clk), .Q(
        \row1_buffer[0][5] ) );
  DFFQXL \row2_buffer_reg[225][4]  ( .D(\row3_buffer[0][4] ), .CK(clk), .Q(
        \row2_buffer[225][4] ) );
  DFFQXL \row2_buffer_reg[224][4]  ( .D(\row2_buffer[225][4] ), .CK(clk), .Q(
        \row2_buffer[224][4] ) );
  DFFQXL \row2_buffer_reg[223][4]  ( .D(\row2_buffer[224][4] ), .CK(clk), .Q(
        \row2_buffer[223][4] ) );
  DFFQXL \row2_buffer_reg[222][4]  ( .D(\row2_buffer[223][4] ), .CK(clk), .Q(
        \row2_buffer[222][4] ) );
  DFFQXL \row2_buffer_reg[221][4]  ( .D(\row2_buffer[222][4] ), .CK(clk), .Q(
        \row2_buffer[221][4] ) );
  DFFQXL \row2_buffer_reg[220][4]  ( .D(\row2_buffer[221][4] ), .CK(clk), .Q(
        \row2_buffer[220][4] ) );
  DFFQXL \row2_buffer_reg[219][4]  ( .D(\row2_buffer[220][4] ), .CK(clk), .Q(
        \row2_buffer[219][4] ) );
  DFFQXL \row2_buffer_reg[218][4]  ( .D(\row2_buffer[219][4] ), .CK(clk), .Q(
        \row2_buffer[218][4] ) );
  DFFQXL \row2_buffer_reg[217][4]  ( .D(\row2_buffer[218][4] ), .CK(clk), .Q(
        \row2_buffer[217][4] ) );
  DFFQXL \row2_buffer_reg[216][4]  ( .D(\row2_buffer[217][4] ), .CK(clk), .Q(
        \row2_buffer[216][4] ) );
  DFFQXL \row2_buffer_reg[215][4]  ( .D(\row2_buffer[216][4] ), .CK(clk), .Q(
        \row2_buffer[215][4] ) );
  DFFQXL \row2_buffer_reg[214][4]  ( .D(\row2_buffer[215][4] ), .CK(clk), .Q(
        \row2_buffer[214][4] ) );
  DFFQXL \row2_buffer_reg[213][4]  ( .D(\row2_buffer[214][4] ), .CK(clk), .Q(
        \row2_buffer[213][4] ) );
  DFFQXL \row2_buffer_reg[212][4]  ( .D(\row2_buffer[213][4] ), .CK(clk), .Q(
        \row2_buffer[212][4] ) );
  DFFQXL \row2_buffer_reg[211][4]  ( .D(\row2_buffer[212][4] ), .CK(clk), .Q(
        \row2_buffer[211][4] ) );
  DFFQXL \row2_buffer_reg[210][4]  ( .D(\row2_buffer[211][4] ), .CK(clk), .Q(
        \row2_buffer[210][4] ) );
  DFFQXL \row2_buffer_reg[209][4]  ( .D(\row2_buffer[210][4] ), .CK(clk), .Q(
        \row2_buffer[209][4] ) );
  DFFQXL \row2_buffer_reg[208][4]  ( .D(\row2_buffer[209][4] ), .CK(clk), .Q(
        \row2_buffer[208][4] ) );
  DFFQXL \row2_buffer_reg[207][4]  ( .D(\row2_buffer[208][4] ), .CK(clk), .Q(
        \row2_buffer[207][4] ) );
  DFFQXL \row2_buffer_reg[206][4]  ( .D(\row2_buffer[207][4] ), .CK(clk), .Q(
        \row2_buffer[206][4] ) );
  DFFQXL \row2_buffer_reg[205][4]  ( .D(\row2_buffer[206][4] ), .CK(clk), .Q(
        \row2_buffer[205][4] ) );
  DFFQXL \row2_buffer_reg[204][4]  ( .D(\row2_buffer[205][4] ), .CK(clk), .Q(
        \row2_buffer[204][4] ) );
  DFFQXL \row2_buffer_reg[203][4]  ( .D(\row2_buffer[204][4] ), .CK(clk), .Q(
        \row2_buffer[203][4] ) );
  DFFQXL \row2_buffer_reg[202][4]  ( .D(\row2_buffer[203][4] ), .CK(clk), .Q(
        \row2_buffer[202][4] ) );
  DFFQXL \row2_buffer_reg[201][4]  ( .D(\row2_buffer[202][4] ), .CK(clk), .Q(
        \row2_buffer[201][4] ) );
  DFFQXL \row2_buffer_reg[200][4]  ( .D(\row2_buffer[201][4] ), .CK(clk), .Q(
        \row2_buffer[200][4] ) );
  DFFQXL \row2_buffer_reg[199][4]  ( .D(\row2_buffer[200][4] ), .CK(clk), .Q(
        \row2_buffer[199][4] ) );
  DFFQXL \row2_buffer_reg[198][4]  ( .D(\row2_buffer[199][4] ), .CK(clk), .Q(
        \row2_buffer[198][4] ) );
  DFFQXL \row2_buffer_reg[197][4]  ( .D(\row2_buffer[198][4] ), .CK(clk), .Q(
        \row2_buffer[197][4] ) );
  DFFQXL \row2_buffer_reg[196][4]  ( .D(\row2_buffer[197][4] ), .CK(clk), .Q(
        \row2_buffer[196][4] ) );
  DFFQXL \row2_buffer_reg[195][4]  ( .D(\row2_buffer[196][4] ), .CK(clk), .Q(
        \row2_buffer[195][4] ) );
  DFFQXL \row2_buffer_reg[194][4]  ( .D(\row2_buffer[195][4] ), .CK(clk), .Q(
        \row2_buffer[194][4] ) );
  DFFQXL \row2_buffer_reg[193][4]  ( .D(\row2_buffer[194][4] ), .CK(clk), .Q(
        \row2_buffer[193][4] ) );
  DFFQXL \row2_buffer_reg[192][4]  ( .D(\row2_buffer[193][4] ), .CK(clk), .Q(
        \row2_buffer[192][4] ) );
  DFFQXL \row2_buffer_reg[191][4]  ( .D(\row2_buffer[192][4] ), .CK(clk), .Q(
        \row2_buffer[191][4] ) );
  DFFQXL \row2_buffer_reg[190][4]  ( .D(\row2_buffer[191][4] ), .CK(clk), .Q(
        \row2_buffer[190][4] ) );
  DFFQXL \row2_buffer_reg[189][4]  ( .D(\row2_buffer[190][4] ), .CK(clk), .Q(
        \row2_buffer[189][4] ) );
  DFFQXL \row2_buffer_reg[188][4]  ( .D(\row2_buffer[189][4] ), .CK(clk), .Q(
        \row2_buffer[188][4] ) );
  DFFQXL \row2_buffer_reg[187][4]  ( .D(\row2_buffer[188][4] ), .CK(clk), .Q(
        \row2_buffer[187][4] ) );
  DFFQXL \row2_buffer_reg[186][4]  ( .D(\row2_buffer[187][4] ), .CK(clk), .Q(
        \row2_buffer[186][4] ) );
  DFFQXL \row2_buffer_reg[185][4]  ( .D(\row2_buffer[186][4] ), .CK(clk), .Q(
        \row2_buffer[185][4] ) );
  DFFQXL \row2_buffer_reg[184][4]  ( .D(\row2_buffer[185][4] ), .CK(clk), .Q(
        \row2_buffer[184][4] ) );
  DFFQXL \row2_buffer_reg[183][4]  ( .D(\row2_buffer[184][4] ), .CK(clk), .Q(
        \row2_buffer[183][4] ) );
  DFFQXL \row2_buffer_reg[182][4]  ( .D(\row2_buffer[183][4] ), .CK(clk), .Q(
        \row2_buffer[182][4] ) );
  DFFQXL \row2_buffer_reg[181][4]  ( .D(\row2_buffer[182][4] ), .CK(clk), .Q(
        \row2_buffer[181][4] ) );
  DFFQXL \row2_buffer_reg[180][4]  ( .D(\row2_buffer[181][4] ), .CK(clk), .Q(
        \row2_buffer[180][4] ) );
  DFFQXL \row2_buffer_reg[179][4]  ( .D(\row2_buffer[180][4] ), .CK(clk), .Q(
        \row2_buffer[179][4] ) );
  DFFQXL \row2_buffer_reg[178][4]  ( .D(\row2_buffer[179][4] ), .CK(clk), .Q(
        \row2_buffer[178][4] ) );
  DFFQXL \row2_buffer_reg[177][4]  ( .D(\row2_buffer[178][4] ), .CK(clk), .Q(
        \row2_buffer[177][4] ) );
  DFFQXL \row2_buffer_reg[176][4]  ( .D(\row2_buffer[177][4] ), .CK(clk), .Q(
        \row2_buffer[176][4] ) );
  DFFQXL \row2_buffer_reg[175][4]  ( .D(\row2_buffer[176][4] ), .CK(clk), .Q(
        \row2_buffer[175][4] ) );
  DFFQXL \row2_buffer_reg[174][4]  ( .D(\row2_buffer[175][4] ), .CK(clk), .Q(
        \row2_buffer[174][4] ) );
  DFFQXL \row2_buffer_reg[173][4]  ( .D(\row2_buffer[174][4] ), .CK(clk), .Q(
        \row2_buffer[173][4] ) );
  DFFQXL \row2_buffer_reg[172][4]  ( .D(\row2_buffer[173][4] ), .CK(clk), .Q(
        \row2_buffer[172][4] ) );
  DFFQXL \row2_buffer_reg[171][4]  ( .D(\row2_buffer[172][4] ), .CK(clk), .Q(
        \row2_buffer[171][4] ) );
  DFFQXL \row2_buffer_reg[170][4]  ( .D(\row2_buffer[171][4] ), .CK(clk), .Q(
        \row2_buffer[170][4] ) );
  DFFQXL \row2_buffer_reg[169][4]  ( .D(\row2_buffer[170][4] ), .CK(clk), .Q(
        \row2_buffer[169][4] ) );
  DFFQXL \row2_buffer_reg[168][4]  ( .D(\row2_buffer[169][4] ), .CK(clk), .Q(
        \row2_buffer[168][4] ) );
  DFFQXL \row2_buffer_reg[167][4]  ( .D(\row2_buffer[168][4] ), .CK(clk), .Q(
        \row2_buffer[167][4] ) );
  DFFQXL \row2_buffer_reg[166][4]  ( .D(\row2_buffer[167][4] ), .CK(clk), .Q(
        \row2_buffer[166][4] ) );
  DFFQXL \row2_buffer_reg[165][4]  ( .D(\row2_buffer[166][4] ), .CK(clk), .Q(
        \row2_buffer[165][4] ) );
  DFFQXL \row2_buffer_reg[164][4]  ( .D(\row2_buffer[165][4] ), .CK(clk), .Q(
        \row2_buffer[164][4] ) );
  DFFQXL \row2_buffer_reg[163][4]  ( .D(\row2_buffer[164][4] ), .CK(clk), .Q(
        \row2_buffer[163][4] ) );
  DFFQXL \row2_buffer_reg[162][4]  ( .D(\row2_buffer[163][4] ), .CK(clk), .Q(
        \row2_buffer[162][4] ) );
  DFFQXL \row2_buffer_reg[161][4]  ( .D(\row2_buffer[162][4] ), .CK(clk), .Q(
        \row2_buffer[161][4] ) );
  DFFQXL \row2_buffer_reg[160][4]  ( .D(\row2_buffer[161][4] ), .CK(clk), .Q(
        \row2_buffer[160][4] ) );
  DFFQXL \row2_buffer_reg[159][4]  ( .D(\row2_buffer[160][4] ), .CK(clk), .Q(
        \row2_buffer[159][4] ) );
  DFFQXL \row2_buffer_reg[158][4]  ( .D(\row2_buffer[159][4] ), .CK(clk), .Q(
        \row2_buffer[158][4] ) );
  DFFQXL \row2_buffer_reg[157][4]  ( .D(\row2_buffer[158][4] ), .CK(clk), .Q(
        \row2_buffer[157][4] ) );
  DFFQXL \row2_buffer_reg[156][4]  ( .D(\row2_buffer[157][4] ), .CK(clk), .Q(
        \row2_buffer[156][4] ) );
  DFFQXL \row2_buffer_reg[155][4]  ( .D(\row2_buffer[156][4] ), .CK(clk), .Q(
        \row2_buffer[155][4] ) );
  DFFQXL \row2_buffer_reg[154][4]  ( .D(\row2_buffer[155][4] ), .CK(clk), .Q(
        \row2_buffer[154][4] ) );
  DFFQXL \row2_buffer_reg[153][4]  ( .D(\row2_buffer[154][4] ), .CK(clk), .Q(
        \row2_buffer[153][4] ) );
  DFFQXL \row2_buffer_reg[152][4]  ( .D(\row2_buffer[153][4] ), .CK(clk), .Q(
        \row2_buffer[152][4] ) );
  DFFQXL \row2_buffer_reg[151][4]  ( .D(\row2_buffer[152][4] ), .CK(clk), .Q(
        \row2_buffer[151][4] ) );
  DFFQXL \row2_buffer_reg[150][4]  ( .D(\row2_buffer[151][4] ), .CK(clk), .Q(
        \row2_buffer[150][4] ) );
  DFFQXL \row2_buffer_reg[149][4]  ( .D(\row2_buffer[150][4] ), .CK(clk), .Q(
        \row2_buffer[149][4] ) );
  DFFQXL \row2_buffer_reg[148][4]  ( .D(\row2_buffer[149][4] ), .CK(clk), .Q(
        \row2_buffer[148][4] ) );
  DFFQXL \row2_buffer_reg[147][4]  ( .D(\row2_buffer[148][4] ), .CK(clk), .Q(
        \row2_buffer[147][4] ) );
  DFFQXL \row2_buffer_reg[146][4]  ( .D(\row2_buffer[147][4] ), .CK(clk), .Q(
        \row2_buffer[146][4] ) );
  DFFQXL \row2_buffer_reg[145][4]  ( .D(\row2_buffer[146][4] ), .CK(clk), .Q(
        \row2_buffer[145][4] ) );
  DFFQXL \row2_buffer_reg[144][4]  ( .D(\row2_buffer[145][4] ), .CK(clk), .Q(
        \row2_buffer[144][4] ) );
  DFFQXL \row2_buffer_reg[143][4]  ( .D(\row2_buffer[144][4] ), .CK(clk), .Q(
        \row2_buffer[143][4] ) );
  DFFQXL \row2_buffer_reg[142][4]  ( .D(\row2_buffer[143][4] ), .CK(clk), .Q(
        \row2_buffer[142][4] ) );
  DFFQXL \row2_buffer_reg[141][4]  ( .D(\row2_buffer[142][4] ), .CK(clk), .Q(
        \row2_buffer[141][4] ) );
  DFFQXL \row2_buffer_reg[140][4]  ( .D(\row2_buffer[141][4] ), .CK(clk), .Q(
        \row2_buffer[140][4] ) );
  DFFQXL \row2_buffer_reg[139][4]  ( .D(\row2_buffer[140][4] ), .CK(clk), .Q(
        \row2_buffer[139][4] ) );
  DFFQXL \row2_buffer_reg[138][4]  ( .D(\row2_buffer[139][4] ), .CK(clk), .Q(
        \row2_buffer[138][4] ) );
  DFFQXL \row2_buffer_reg[137][4]  ( .D(\row2_buffer[138][4] ), .CK(clk), .Q(
        \row2_buffer[137][4] ) );
  DFFQXL \row2_buffer_reg[136][4]  ( .D(\row2_buffer[137][4] ), .CK(clk), .Q(
        \row2_buffer[136][4] ) );
  DFFQXL \row2_buffer_reg[135][4]  ( .D(\row2_buffer[136][4] ), .CK(clk), .Q(
        \row2_buffer[135][4] ) );
  DFFQXL \row2_buffer_reg[134][4]  ( .D(\row2_buffer[135][4] ), .CK(clk), .Q(
        \row2_buffer[134][4] ) );
  DFFQXL \row2_buffer_reg[133][4]  ( .D(\row2_buffer[134][4] ), .CK(clk), .Q(
        \row2_buffer[133][4] ) );
  DFFQXL \row2_buffer_reg[132][4]  ( .D(\row2_buffer[133][4] ), .CK(clk), .Q(
        \row2_buffer[132][4] ) );
  DFFQXL \row2_buffer_reg[131][4]  ( .D(\row2_buffer[132][4] ), .CK(clk), .Q(
        \row2_buffer[131][4] ) );
  DFFQXL \row2_buffer_reg[130][4]  ( .D(\row2_buffer[131][4] ), .CK(clk), .Q(
        \row2_buffer[130][4] ) );
  DFFQXL \row2_buffer_reg[129][4]  ( .D(\row2_buffer[130][4] ), .CK(clk), .Q(
        \row2_buffer[129][4] ) );
  DFFQXL \row2_buffer_reg[128][4]  ( .D(\row2_buffer[129][4] ), .CK(clk), .Q(
        \row2_buffer[128][4] ) );
  DFFQXL \row2_buffer_reg[127][4]  ( .D(\row2_buffer[128][4] ), .CK(clk), .Q(
        \row2_buffer[127][4] ) );
  DFFQXL \row2_buffer_reg[126][4]  ( .D(\row2_buffer[127][4] ), .CK(clk), .Q(
        \row2_buffer[126][4] ) );
  DFFQXL \row2_buffer_reg[125][4]  ( .D(\row2_buffer[126][4] ), .CK(clk), .Q(
        \row2_buffer[125][4] ) );
  DFFQXL \row2_buffer_reg[124][4]  ( .D(\row2_buffer[125][4] ), .CK(clk), .Q(
        \row2_buffer[124][4] ) );
  DFFQXL \row2_buffer_reg[123][4]  ( .D(\row2_buffer[124][4] ), .CK(clk), .Q(
        \row2_buffer[123][4] ) );
  DFFQXL \row2_buffer_reg[122][4]  ( .D(\row2_buffer[123][4] ), .CK(clk), .Q(
        \row2_buffer[122][4] ) );
  DFFQXL \row2_buffer_reg[121][4]  ( .D(\row2_buffer[122][4] ), .CK(clk), .Q(
        \row2_buffer[121][4] ) );
  DFFQXL \row2_buffer_reg[120][4]  ( .D(\row2_buffer[121][4] ), .CK(clk), .Q(
        \row2_buffer[120][4] ) );
  DFFQXL \row2_buffer_reg[119][4]  ( .D(\row2_buffer[120][4] ), .CK(clk), .Q(
        \row2_buffer[119][4] ) );
  DFFQXL \row2_buffer_reg[118][4]  ( .D(\row2_buffer[119][4] ), .CK(clk), .Q(
        \row2_buffer[118][4] ) );
  DFFQXL \row2_buffer_reg[117][4]  ( .D(\row2_buffer[118][4] ), .CK(clk), .Q(
        \row2_buffer[117][4] ) );
  DFFQXL \row2_buffer_reg[116][4]  ( .D(\row2_buffer[117][4] ), .CK(clk), .Q(
        \row2_buffer[116][4] ) );
  DFFQXL \row2_buffer_reg[115][4]  ( .D(\row2_buffer[116][4] ), .CK(clk), .Q(
        \row2_buffer[115][4] ) );
  DFFQXL \row2_buffer_reg[114][4]  ( .D(\row2_buffer[115][4] ), .CK(clk), .Q(
        \row2_buffer[114][4] ) );
  DFFQXL \row2_buffer_reg[113][4]  ( .D(\row2_buffer[114][4] ), .CK(clk), .Q(
        \row2_buffer[113][4] ) );
  DFFQXL \row2_buffer_reg[112][4]  ( .D(\row2_buffer[113][4] ), .CK(clk), .Q(
        \row2_buffer[112][4] ) );
  DFFQXL \row2_buffer_reg[111][4]  ( .D(\row2_buffer[112][4] ), .CK(clk), .Q(
        \row2_buffer[111][4] ) );
  DFFQXL \row2_buffer_reg[110][4]  ( .D(\row2_buffer[111][4] ), .CK(clk), .Q(
        \row2_buffer[110][4] ) );
  DFFQXL \row2_buffer_reg[109][4]  ( .D(\row2_buffer[110][4] ), .CK(clk), .Q(
        \row2_buffer[109][4] ) );
  DFFQXL \row2_buffer_reg[108][4]  ( .D(\row2_buffer[109][4] ), .CK(clk), .Q(
        \row2_buffer[108][4] ) );
  DFFQXL \row2_buffer_reg[107][4]  ( .D(\row2_buffer[108][4] ), .CK(clk), .Q(
        \row2_buffer[107][4] ) );
  DFFQXL \row2_buffer_reg[106][4]  ( .D(\row2_buffer[107][4] ), .CK(clk), .Q(
        \row2_buffer[106][4] ) );
  DFFQXL \row2_buffer_reg[105][4]  ( .D(\row2_buffer[106][4] ), .CK(clk), .Q(
        \row2_buffer[105][4] ) );
  DFFQXL \row2_buffer_reg[104][4]  ( .D(\row2_buffer[105][4] ), .CK(clk), .Q(
        \row2_buffer[104][4] ) );
  DFFQXL \row2_buffer_reg[103][4]  ( .D(\row2_buffer[104][4] ), .CK(clk), .Q(
        \row2_buffer[103][4] ) );
  DFFQXL \row2_buffer_reg[102][4]  ( .D(\row2_buffer[103][4] ), .CK(clk), .Q(
        \row2_buffer[102][4] ) );
  DFFQXL \row2_buffer_reg[101][4]  ( .D(\row2_buffer[102][4] ), .CK(clk), .Q(
        \row2_buffer[101][4] ) );
  DFFQXL \row2_buffer_reg[100][4]  ( .D(\row2_buffer[101][4] ), .CK(clk), .Q(
        \row2_buffer[100][4] ) );
  DFFQXL \row2_buffer_reg[99][4]  ( .D(\row2_buffer[100][4] ), .CK(clk), .Q(
        \row2_buffer[99][4] ) );
  DFFQXL \row2_buffer_reg[98][4]  ( .D(\row2_buffer[99][4] ), .CK(clk), .Q(
        \row2_buffer[98][4] ) );
  DFFQXL \row2_buffer_reg[97][4]  ( .D(\row2_buffer[98][4] ), .CK(clk), .Q(
        \row2_buffer[97][4] ) );
  DFFQXL \row2_buffer_reg[96][4]  ( .D(\row2_buffer[97][4] ), .CK(clk), .Q(
        \row2_buffer[96][4] ) );
  DFFQXL \row2_buffer_reg[95][4]  ( .D(\row2_buffer[96][4] ), .CK(clk), .Q(
        \row2_buffer[95][4] ) );
  DFFQXL \row2_buffer_reg[94][4]  ( .D(\row2_buffer[95][4] ), .CK(clk), .Q(
        \row2_buffer[94][4] ) );
  DFFQXL \row2_buffer_reg[93][4]  ( .D(\row2_buffer[94][4] ), .CK(clk), .Q(
        \row2_buffer[93][4] ) );
  DFFQXL \row2_buffer_reg[92][4]  ( .D(\row2_buffer[93][4] ), .CK(clk), .Q(
        \row2_buffer[92][4] ) );
  DFFQXL \row2_buffer_reg[91][4]  ( .D(\row2_buffer[92][4] ), .CK(clk), .Q(
        \row2_buffer[91][4] ) );
  DFFQXL \row2_buffer_reg[90][4]  ( .D(\row2_buffer[91][4] ), .CK(clk), .Q(
        \row2_buffer[90][4] ) );
  DFFQXL \row2_buffer_reg[89][4]  ( .D(\row2_buffer[90][4] ), .CK(clk), .Q(
        \row2_buffer[89][4] ) );
  DFFQXL \row2_buffer_reg[88][4]  ( .D(\row2_buffer[89][4] ), .CK(clk), .Q(
        \row2_buffer[88][4] ) );
  DFFQXL \row2_buffer_reg[87][4]  ( .D(\row2_buffer[88][4] ), .CK(clk), .Q(
        \row2_buffer[87][4] ) );
  DFFQXL \row2_buffer_reg[86][4]  ( .D(\row2_buffer[87][4] ), .CK(clk), .Q(
        \row2_buffer[86][4] ) );
  DFFQXL \row2_buffer_reg[85][4]  ( .D(\row2_buffer[86][4] ), .CK(clk), .Q(
        \row2_buffer[85][4] ) );
  DFFQXL \row2_buffer_reg[84][4]  ( .D(\row2_buffer[85][4] ), .CK(clk), .Q(
        \row2_buffer[84][4] ) );
  DFFQXL \row2_buffer_reg[83][4]  ( .D(\row2_buffer[84][4] ), .CK(clk), .Q(
        \row2_buffer[83][4] ) );
  DFFQXL \row2_buffer_reg[82][4]  ( .D(\row2_buffer[83][4] ), .CK(clk), .Q(
        \row2_buffer[82][4] ) );
  DFFQXL \row2_buffer_reg[81][4]  ( .D(\row2_buffer[82][4] ), .CK(clk), .Q(
        \row2_buffer[81][4] ) );
  DFFQXL \row2_buffer_reg[80][4]  ( .D(\row2_buffer[81][4] ), .CK(clk), .Q(
        \row2_buffer[80][4] ) );
  DFFQXL \row2_buffer_reg[79][4]  ( .D(\row2_buffer[80][4] ), .CK(clk), .Q(
        \row2_buffer[79][4] ) );
  DFFQXL \row2_buffer_reg[78][4]  ( .D(\row2_buffer[79][4] ), .CK(clk), .Q(
        \row2_buffer[78][4] ) );
  DFFQXL \row2_buffer_reg[77][4]  ( .D(\row2_buffer[78][4] ), .CK(clk), .Q(
        \row2_buffer[77][4] ) );
  DFFQXL \row2_buffer_reg[76][4]  ( .D(\row2_buffer[77][4] ), .CK(clk), .Q(
        \row2_buffer[76][4] ) );
  DFFQXL \row2_buffer_reg[75][4]  ( .D(\row2_buffer[76][4] ), .CK(clk), .Q(
        \row2_buffer[75][4] ) );
  DFFQXL \row2_buffer_reg[74][4]  ( .D(\row2_buffer[75][4] ), .CK(clk), .Q(
        \row2_buffer[74][4] ) );
  DFFQXL \row2_buffer_reg[73][4]  ( .D(\row2_buffer[74][4] ), .CK(clk), .Q(
        \row2_buffer[73][4] ) );
  DFFQXL \row2_buffer_reg[72][4]  ( .D(\row2_buffer[73][4] ), .CK(clk), .Q(
        \row2_buffer[72][4] ) );
  DFFQXL \row2_buffer_reg[71][4]  ( .D(\row2_buffer[72][4] ), .CK(clk), .Q(
        \row2_buffer[71][4] ) );
  DFFQXL \row2_buffer_reg[70][4]  ( .D(\row2_buffer[71][4] ), .CK(clk), .Q(
        \row2_buffer[70][4] ) );
  DFFQXL \row2_buffer_reg[69][4]  ( .D(\row2_buffer[70][4] ), .CK(clk), .Q(
        \row2_buffer[69][4] ) );
  DFFQXL \row2_buffer_reg[68][4]  ( .D(\row2_buffer[69][4] ), .CK(clk), .Q(
        \row2_buffer[68][4] ) );
  DFFQXL \row2_buffer_reg[67][4]  ( .D(\row2_buffer[68][4] ), .CK(clk), .Q(
        \row2_buffer[67][4] ) );
  DFFQXL \row2_buffer_reg[66][4]  ( .D(\row2_buffer[67][4] ), .CK(clk), .Q(
        \row2_buffer[66][4] ) );
  DFFQXL \row2_buffer_reg[65][4]  ( .D(\row2_buffer[66][4] ), .CK(clk), .Q(
        \row2_buffer[65][4] ) );
  DFFQXL \row2_buffer_reg[64][4]  ( .D(\row2_buffer[65][4] ), .CK(clk), .Q(
        \row2_buffer[64][4] ) );
  DFFQXL \row2_buffer_reg[63][4]  ( .D(\row2_buffer[64][4] ), .CK(clk), .Q(
        \row2_buffer[63][4] ) );
  DFFQXL \row2_buffer_reg[62][4]  ( .D(\row2_buffer[63][4] ), .CK(clk), .Q(
        \row2_buffer[62][4] ) );
  DFFQXL \row2_buffer_reg[61][4]  ( .D(\row2_buffer[62][4] ), .CK(clk), .Q(
        \row2_buffer[61][4] ) );
  DFFQXL \row2_buffer_reg[60][4]  ( .D(\row2_buffer[61][4] ), .CK(clk), .Q(
        \row2_buffer[60][4] ) );
  DFFQXL \row2_buffer_reg[59][4]  ( .D(\row2_buffer[60][4] ), .CK(clk), .Q(
        \row2_buffer[59][4] ) );
  DFFQXL \row2_buffer_reg[58][4]  ( .D(\row2_buffer[59][4] ), .CK(clk), .Q(
        \row2_buffer[58][4] ) );
  DFFQXL \row2_buffer_reg[57][4]  ( .D(\row2_buffer[58][4] ), .CK(clk), .Q(
        \row2_buffer[57][4] ) );
  DFFQXL \row2_buffer_reg[56][4]  ( .D(\row2_buffer[57][4] ), .CK(clk), .Q(
        \row2_buffer[56][4] ) );
  DFFQXL \row2_buffer_reg[55][4]  ( .D(\row2_buffer[56][4] ), .CK(clk), .Q(
        \row2_buffer[55][4] ) );
  DFFQXL \row2_buffer_reg[54][4]  ( .D(\row2_buffer[55][4] ), .CK(clk), .Q(
        \row2_buffer[54][4] ) );
  DFFQXL \row2_buffer_reg[53][4]  ( .D(\row2_buffer[54][4] ), .CK(clk), .Q(
        \row2_buffer[53][4] ) );
  DFFQXL \row2_buffer_reg[52][4]  ( .D(\row2_buffer[53][4] ), .CK(clk), .Q(
        \row2_buffer[52][4] ) );
  DFFQXL \row2_buffer_reg[51][4]  ( .D(\row2_buffer[52][4] ), .CK(clk), .Q(
        \row2_buffer[51][4] ) );
  DFFQXL \row2_buffer_reg[50][4]  ( .D(\row2_buffer[51][4] ), .CK(clk), .Q(
        \row2_buffer[50][4] ) );
  DFFQXL \row2_buffer_reg[49][4]  ( .D(\row2_buffer[50][4] ), .CK(clk), .Q(
        \row2_buffer[49][4] ) );
  DFFQXL \row2_buffer_reg[48][4]  ( .D(\row2_buffer[49][4] ), .CK(clk), .Q(
        \row2_buffer[48][4] ) );
  DFFQXL \row2_buffer_reg[47][4]  ( .D(\row2_buffer[48][4] ), .CK(clk), .Q(
        \row2_buffer[47][4] ) );
  DFFQXL \row2_buffer_reg[46][4]  ( .D(\row2_buffer[47][4] ), .CK(clk), .Q(
        \row2_buffer[46][4] ) );
  DFFQXL \row2_buffer_reg[45][4]  ( .D(\row2_buffer[46][4] ), .CK(clk), .Q(
        \row2_buffer[45][4] ) );
  DFFQXL \row2_buffer_reg[44][4]  ( .D(\row2_buffer[45][4] ), .CK(clk), .Q(
        \row2_buffer[44][4] ) );
  DFFQXL \row2_buffer_reg[43][4]  ( .D(\row2_buffer[44][4] ), .CK(clk), .Q(
        \row2_buffer[43][4] ) );
  DFFQXL \row2_buffer_reg[42][4]  ( .D(\row2_buffer[43][4] ), .CK(clk), .Q(
        \row2_buffer[42][4] ) );
  DFFQXL \row2_buffer_reg[41][4]  ( .D(\row2_buffer[42][4] ), .CK(clk), .Q(
        \row2_buffer[41][4] ) );
  DFFQXL \row2_buffer_reg[40][4]  ( .D(\row2_buffer[41][4] ), .CK(clk), .Q(
        \row2_buffer[40][4] ) );
  DFFQXL \row2_buffer_reg[39][4]  ( .D(\row2_buffer[40][4] ), .CK(clk), .Q(
        \row2_buffer[39][4] ) );
  DFFQXL \row2_buffer_reg[38][4]  ( .D(\row2_buffer[39][4] ), .CK(clk), .Q(
        \row2_buffer[38][4] ) );
  DFFQXL \row2_buffer_reg[37][4]  ( .D(\row2_buffer[38][4] ), .CK(clk), .Q(
        \row2_buffer[37][4] ) );
  DFFQXL \row2_buffer_reg[36][4]  ( .D(\row2_buffer[37][4] ), .CK(clk), .Q(
        \row2_buffer[36][4] ) );
  DFFQXL \row2_buffer_reg[35][4]  ( .D(\row2_buffer[36][4] ), .CK(clk), .Q(
        \row2_buffer[35][4] ) );
  DFFQXL \row2_buffer_reg[34][4]  ( .D(\row2_buffer[35][4] ), .CK(clk), .Q(
        \row2_buffer[34][4] ) );
  DFFQXL \row2_buffer_reg[33][4]  ( .D(\row2_buffer[34][4] ), .CK(clk), .Q(
        \row2_buffer[33][4] ) );
  DFFQXL \row2_buffer_reg[32][4]  ( .D(\row2_buffer[33][4] ), .CK(clk), .Q(
        \row2_buffer[32][4] ) );
  DFFQXL \row2_buffer_reg[31][4]  ( .D(\row2_buffer[32][4] ), .CK(clk), .Q(
        \row2_buffer[31][4] ) );
  DFFQXL \row2_buffer_reg[30][4]  ( .D(\row2_buffer[31][4] ), .CK(clk), .Q(
        \row2_buffer[30][4] ) );
  DFFQXL \row2_buffer_reg[29][4]  ( .D(\row2_buffer[30][4] ), .CK(clk), .Q(
        \row2_buffer[29][4] ) );
  DFFQXL \row2_buffer_reg[28][4]  ( .D(\row2_buffer[29][4] ), .CK(clk), .Q(
        \row2_buffer[28][4] ) );
  DFFQXL \row2_buffer_reg[27][4]  ( .D(\row2_buffer[28][4] ), .CK(clk), .Q(
        \row2_buffer[27][4] ) );
  DFFQXL \row2_buffer_reg[26][4]  ( .D(\row2_buffer[27][4] ), .CK(clk), .Q(
        \row2_buffer[26][4] ) );
  DFFQXL \row2_buffer_reg[25][4]  ( .D(\row2_buffer[26][4] ), .CK(clk), .Q(
        \row2_buffer[25][4] ) );
  DFFQXL \row2_buffer_reg[24][4]  ( .D(\row2_buffer[25][4] ), .CK(clk), .Q(
        \row2_buffer[24][4] ) );
  DFFQXL \row2_buffer_reg[23][4]  ( .D(\row2_buffer[24][4] ), .CK(clk), .Q(
        \row2_buffer[23][4] ) );
  DFFQXL \row2_buffer_reg[22][4]  ( .D(\row2_buffer[23][4] ), .CK(clk), .Q(
        \row2_buffer[22][4] ) );
  DFFQXL \row2_buffer_reg[21][4]  ( .D(\row2_buffer[22][4] ), .CK(clk), .Q(
        \row2_buffer[21][4] ) );
  DFFQXL \row2_buffer_reg[20][4]  ( .D(\row2_buffer[21][4] ), .CK(clk), .Q(
        \row2_buffer[20][4] ) );
  DFFQXL \row2_buffer_reg[19][4]  ( .D(\row2_buffer[20][4] ), .CK(clk), .Q(
        \row2_buffer[19][4] ) );
  DFFQXL \row2_buffer_reg[18][4]  ( .D(\row2_buffer[19][4] ), .CK(clk), .Q(
        \row2_buffer[18][4] ) );
  DFFQXL \row2_buffer_reg[17][4]  ( .D(\row2_buffer[18][4] ), .CK(clk), .Q(
        \row2_buffer[17][4] ) );
  DFFQXL \row2_buffer_reg[16][4]  ( .D(\row2_buffer[17][4] ), .CK(clk), .Q(
        \row2_buffer[16][4] ) );
  DFFQXL \row2_buffer_reg[15][4]  ( .D(\row2_buffer[16][4] ), .CK(clk), .Q(
        \row2_buffer[15][4] ) );
  DFFQXL \row2_buffer_reg[14][4]  ( .D(\row2_buffer[15][4] ), .CK(clk), .Q(
        \row2_buffer[14][4] ) );
  DFFQXL \row2_buffer_reg[13][4]  ( .D(\row2_buffer[14][4] ), .CK(clk), .Q(
        \row2_buffer[13][4] ) );
  DFFQXL \row2_buffer_reg[12][4]  ( .D(\row2_buffer[13][4] ), .CK(clk), .Q(
        \row2_buffer[12][4] ) );
  DFFQXL \row2_buffer_reg[11][4]  ( .D(\row2_buffer[12][4] ), .CK(clk), .Q(
        \row2_buffer[11][4] ) );
  DFFQXL \row2_buffer_reg[10][4]  ( .D(\row2_buffer[11][4] ), .CK(clk), .Q(
        \row2_buffer[10][4] ) );
  DFFQXL \row2_buffer_reg[9][4]  ( .D(\row2_buffer[10][4] ), .CK(clk), .Q(
        \row2_buffer[9][4] ) );
  DFFQXL \row2_buffer_reg[8][4]  ( .D(\row2_buffer[9][4] ), .CK(clk), .Q(
        \row2_buffer[8][4] ) );
  DFFQXL \row2_buffer_reg[7][4]  ( .D(\row2_buffer[8][4] ), .CK(clk), .Q(
        \row2_buffer[7][4] ) );
  DFFQXL \row2_buffer_reg[6][4]  ( .D(\row2_buffer[7][4] ), .CK(clk), .Q(
        \row2_buffer[6][4] ) );
  DFFQXL \row2_buffer_reg[5][4]  ( .D(\row2_buffer[6][4] ), .CK(clk), .Q(
        \row2_buffer[5][4] ) );
  DFFQXL \row2_buffer_reg[4][4]  ( .D(\row2_buffer[5][4] ), .CK(clk), .Q(
        \row2_buffer[4][4] ) );
  DFFQXL \row2_buffer_reg[3][4]  ( .D(\row2_buffer[4][4] ), .CK(clk), .Q(
        \row2_buffer[3][4] ) );
  DFFQXL \row1_buffer_reg[225][4]  ( .D(\row2_buffer[0][4] ), .CK(clk), .Q(
        \row1_buffer[225][4] ) );
  DFFQXL \row1_buffer_reg[224][4]  ( .D(\row1_buffer[225][4] ), .CK(clk), .Q(
        \row1_buffer[224][4] ) );
  DFFQXL \row1_buffer_reg[223][4]  ( .D(\row1_buffer[224][4] ), .CK(clk), .Q(
        \row1_buffer[223][4] ) );
  DFFQXL \row1_buffer_reg[222][4]  ( .D(\row1_buffer[223][4] ), .CK(clk), .Q(
        \row1_buffer[222][4] ) );
  DFFQXL \row1_buffer_reg[221][4]  ( .D(\row1_buffer[222][4] ), .CK(clk), .Q(
        \row1_buffer[221][4] ) );
  DFFQXL \row1_buffer_reg[220][4]  ( .D(\row1_buffer[221][4] ), .CK(clk), .Q(
        \row1_buffer[220][4] ) );
  DFFQXL \row1_buffer_reg[219][4]  ( .D(\row1_buffer[220][4] ), .CK(clk), .Q(
        \row1_buffer[219][4] ) );
  DFFQXL \row1_buffer_reg[218][4]  ( .D(\row1_buffer[219][4] ), .CK(clk), .Q(
        \row1_buffer[218][4] ) );
  DFFQXL \row1_buffer_reg[217][4]  ( .D(\row1_buffer[218][4] ), .CK(clk), .Q(
        \row1_buffer[217][4] ) );
  DFFQXL \row1_buffer_reg[216][4]  ( .D(\row1_buffer[217][4] ), .CK(clk), .Q(
        \row1_buffer[216][4] ) );
  DFFQXL \row1_buffer_reg[215][4]  ( .D(\row1_buffer[216][4] ), .CK(clk), .Q(
        \row1_buffer[215][4] ) );
  DFFQXL \row1_buffer_reg[214][4]  ( .D(\row1_buffer[215][4] ), .CK(clk), .Q(
        \row1_buffer[214][4] ) );
  DFFQXL \row1_buffer_reg[213][4]  ( .D(\row1_buffer[214][4] ), .CK(clk), .Q(
        \row1_buffer[213][4] ) );
  DFFQXL \row1_buffer_reg[212][4]  ( .D(\row1_buffer[213][4] ), .CK(clk), .Q(
        \row1_buffer[212][4] ) );
  DFFQXL \row1_buffer_reg[211][4]  ( .D(\row1_buffer[212][4] ), .CK(clk), .Q(
        \row1_buffer[211][4] ) );
  DFFQXL \row1_buffer_reg[210][4]  ( .D(\row1_buffer[211][4] ), .CK(clk), .Q(
        \row1_buffer[210][4] ) );
  DFFQXL \row1_buffer_reg[209][4]  ( .D(\row1_buffer[210][4] ), .CK(clk), .Q(
        \row1_buffer[209][4] ) );
  DFFQXL \row1_buffer_reg[208][4]  ( .D(\row1_buffer[209][4] ), .CK(clk), .Q(
        \row1_buffer[208][4] ) );
  DFFQXL \row1_buffer_reg[207][4]  ( .D(\row1_buffer[208][4] ), .CK(clk), .Q(
        \row1_buffer[207][4] ) );
  DFFQXL \row1_buffer_reg[206][4]  ( .D(\row1_buffer[207][4] ), .CK(clk), .Q(
        \row1_buffer[206][4] ) );
  DFFQXL \row1_buffer_reg[205][4]  ( .D(\row1_buffer[206][4] ), .CK(clk), .Q(
        \row1_buffer[205][4] ) );
  DFFQXL \row1_buffer_reg[204][4]  ( .D(\row1_buffer[205][4] ), .CK(clk), .Q(
        \row1_buffer[204][4] ) );
  DFFQXL \row1_buffer_reg[203][4]  ( .D(\row1_buffer[204][4] ), .CK(clk), .Q(
        \row1_buffer[203][4] ) );
  DFFQXL \row1_buffer_reg[202][4]  ( .D(\row1_buffer[203][4] ), .CK(clk), .Q(
        \row1_buffer[202][4] ) );
  DFFQXL \row1_buffer_reg[201][4]  ( .D(\row1_buffer[202][4] ), .CK(clk), .Q(
        \row1_buffer[201][4] ) );
  DFFQXL \row1_buffer_reg[200][4]  ( .D(\row1_buffer[201][4] ), .CK(clk), .Q(
        \row1_buffer[200][4] ) );
  DFFQXL \row1_buffer_reg[199][4]  ( .D(\row1_buffer[200][4] ), .CK(clk), .Q(
        \row1_buffer[199][4] ) );
  DFFQXL \row1_buffer_reg[198][4]  ( .D(\row1_buffer[199][4] ), .CK(clk), .Q(
        \row1_buffer[198][4] ) );
  DFFQXL \row1_buffer_reg[197][4]  ( .D(\row1_buffer[198][4] ), .CK(clk), .Q(
        \row1_buffer[197][4] ) );
  DFFQXL \row1_buffer_reg[196][4]  ( .D(\row1_buffer[197][4] ), .CK(clk), .Q(
        \row1_buffer[196][4] ) );
  DFFQXL \row1_buffer_reg[195][4]  ( .D(\row1_buffer[196][4] ), .CK(clk), .Q(
        \row1_buffer[195][4] ) );
  DFFQXL \row1_buffer_reg[194][4]  ( .D(\row1_buffer[195][4] ), .CK(clk), .Q(
        \row1_buffer[194][4] ) );
  DFFQXL \row1_buffer_reg[193][4]  ( .D(\row1_buffer[194][4] ), .CK(clk), .Q(
        \row1_buffer[193][4] ) );
  DFFQXL \row1_buffer_reg[192][4]  ( .D(\row1_buffer[193][4] ), .CK(clk), .Q(
        \row1_buffer[192][4] ) );
  DFFQXL \row1_buffer_reg[191][4]  ( .D(\row1_buffer[192][4] ), .CK(clk), .Q(
        \row1_buffer[191][4] ) );
  DFFQXL \row1_buffer_reg[190][4]  ( .D(\row1_buffer[191][4] ), .CK(clk), .Q(
        \row1_buffer[190][4] ) );
  DFFQXL \row1_buffer_reg[189][4]  ( .D(\row1_buffer[190][4] ), .CK(clk), .Q(
        \row1_buffer[189][4] ) );
  DFFQXL \row1_buffer_reg[188][4]  ( .D(\row1_buffer[189][4] ), .CK(clk), .Q(
        \row1_buffer[188][4] ) );
  DFFQXL \row1_buffer_reg[187][4]  ( .D(\row1_buffer[188][4] ), .CK(clk), .Q(
        \row1_buffer[187][4] ) );
  DFFQXL \row1_buffer_reg[186][4]  ( .D(\row1_buffer[187][4] ), .CK(clk), .Q(
        \row1_buffer[186][4] ) );
  DFFQXL \row1_buffer_reg[185][4]  ( .D(\row1_buffer[186][4] ), .CK(clk), .Q(
        \row1_buffer[185][4] ) );
  DFFQXL \row1_buffer_reg[184][4]  ( .D(\row1_buffer[185][4] ), .CK(clk), .Q(
        \row1_buffer[184][4] ) );
  DFFQXL \row1_buffer_reg[183][4]  ( .D(\row1_buffer[184][4] ), .CK(clk), .Q(
        \row1_buffer[183][4] ) );
  DFFQXL \row1_buffer_reg[182][4]  ( .D(\row1_buffer[183][4] ), .CK(clk), .Q(
        \row1_buffer[182][4] ) );
  DFFQXL \row1_buffer_reg[181][4]  ( .D(\row1_buffer[182][4] ), .CK(clk), .Q(
        \row1_buffer[181][4] ) );
  DFFQXL \row1_buffer_reg[180][4]  ( .D(\row1_buffer[181][4] ), .CK(clk), .Q(
        \row1_buffer[180][4] ) );
  DFFQXL \row1_buffer_reg[179][4]  ( .D(\row1_buffer[180][4] ), .CK(clk), .Q(
        \row1_buffer[179][4] ) );
  DFFQXL \row1_buffer_reg[178][4]  ( .D(\row1_buffer[179][4] ), .CK(clk), .Q(
        \row1_buffer[178][4] ) );
  DFFQXL \row1_buffer_reg[177][4]  ( .D(\row1_buffer[178][4] ), .CK(clk), .Q(
        \row1_buffer[177][4] ) );
  DFFQXL \row1_buffer_reg[176][4]  ( .D(\row1_buffer[177][4] ), .CK(clk), .Q(
        \row1_buffer[176][4] ) );
  DFFQXL \row1_buffer_reg[175][4]  ( .D(\row1_buffer[176][4] ), .CK(clk), .Q(
        \row1_buffer[175][4] ) );
  DFFQXL \row1_buffer_reg[174][4]  ( .D(\row1_buffer[175][4] ), .CK(clk), .Q(
        \row1_buffer[174][4] ) );
  DFFQXL \row1_buffer_reg[173][4]  ( .D(\row1_buffer[174][4] ), .CK(clk), .Q(
        \row1_buffer[173][4] ) );
  DFFQXL \row1_buffer_reg[172][4]  ( .D(\row1_buffer[173][4] ), .CK(clk), .Q(
        \row1_buffer[172][4] ) );
  DFFQXL \row1_buffer_reg[171][4]  ( .D(\row1_buffer[172][4] ), .CK(clk), .Q(
        \row1_buffer[171][4] ) );
  DFFQXL \row1_buffer_reg[170][4]  ( .D(\row1_buffer[171][4] ), .CK(clk), .Q(
        \row1_buffer[170][4] ) );
  DFFQXL \row1_buffer_reg[169][4]  ( .D(\row1_buffer[170][4] ), .CK(clk), .Q(
        \row1_buffer[169][4] ) );
  DFFQXL \row1_buffer_reg[168][4]  ( .D(\row1_buffer[169][4] ), .CK(clk), .Q(
        \row1_buffer[168][4] ) );
  DFFQXL \row1_buffer_reg[167][4]  ( .D(\row1_buffer[168][4] ), .CK(clk), .Q(
        \row1_buffer[167][4] ) );
  DFFQXL \row1_buffer_reg[166][4]  ( .D(\row1_buffer[167][4] ), .CK(clk), .Q(
        \row1_buffer[166][4] ) );
  DFFQXL \row1_buffer_reg[165][4]  ( .D(\row1_buffer[166][4] ), .CK(clk), .Q(
        \row1_buffer[165][4] ) );
  DFFQXL \row1_buffer_reg[164][4]  ( .D(\row1_buffer[165][4] ), .CK(clk), .Q(
        \row1_buffer[164][4] ) );
  DFFQXL \row1_buffer_reg[163][4]  ( .D(\row1_buffer[164][4] ), .CK(clk), .Q(
        \row1_buffer[163][4] ) );
  DFFQXL \row1_buffer_reg[162][4]  ( .D(\row1_buffer[163][4] ), .CK(clk), .Q(
        \row1_buffer[162][4] ) );
  DFFQXL \row1_buffer_reg[161][4]  ( .D(\row1_buffer[162][4] ), .CK(clk), .Q(
        \row1_buffer[161][4] ) );
  DFFQXL \row1_buffer_reg[160][4]  ( .D(\row1_buffer[161][4] ), .CK(clk), .Q(
        \row1_buffer[160][4] ) );
  DFFQXL \row1_buffer_reg[159][4]  ( .D(\row1_buffer[160][4] ), .CK(clk), .Q(
        \row1_buffer[159][4] ) );
  DFFQXL \row1_buffer_reg[158][4]  ( .D(\row1_buffer[159][4] ), .CK(clk), .Q(
        \row1_buffer[158][4] ) );
  DFFQXL \row1_buffer_reg[157][4]  ( .D(\row1_buffer[158][4] ), .CK(clk), .Q(
        \row1_buffer[157][4] ) );
  DFFQXL \row1_buffer_reg[156][4]  ( .D(\row1_buffer[157][4] ), .CK(clk), .Q(
        \row1_buffer[156][4] ) );
  DFFQXL \row1_buffer_reg[155][4]  ( .D(\row1_buffer[156][4] ), .CK(clk), .Q(
        \row1_buffer[155][4] ) );
  DFFQXL \row1_buffer_reg[154][4]  ( .D(\row1_buffer[155][4] ), .CK(clk), .Q(
        \row1_buffer[154][4] ) );
  DFFQXL \row1_buffer_reg[153][4]  ( .D(\row1_buffer[154][4] ), .CK(clk), .Q(
        \row1_buffer[153][4] ) );
  DFFQXL \row1_buffer_reg[152][4]  ( .D(\row1_buffer[153][4] ), .CK(clk), .Q(
        \row1_buffer[152][4] ) );
  DFFQXL \row1_buffer_reg[151][4]  ( .D(\row1_buffer[152][4] ), .CK(clk), .Q(
        \row1_buffer[151][4] ) );
  DFFQXL \row1_buffer_reg[150][4]  ( .D(\row1_buffer[151][4] ), .CK(clk), .Q(
        \row1_buffer[150][4] ) );
  DFFQXL \row1_buffer_reg[149][4]  ( .D(\row1_buffer[150][4] ), .CK(clk), .Q(
        \row1_buffer[149][4] ) );
  DFFQXL \row1_buffer_reg[148][4]  ( .D(\row1_buffer[149][4] ), .CK(clk), .Q(
        \row1_buffer[148][4] ) );
  DFFQXL \row1_buffer_reg[147][4]  ( .D(\row1_buffer[148][4] ), .CK(clk), .Q(
        \row1_buffer[147][4] ) );
  DFFQXL \row1_buffer_reg[146][4]  ( .D(\row1_buffer[147][4] ), .CK(clk), .Q(
        \row1_buffer[146][4] ) );
  DFFQXL \row1_buffer_reg[145][4]  ( .D(\row1_buffer[146][4] ), .CK(clk), .Q(
        \row1_buffer[145][4] ) );
  DFFQXL \row1_buffer_reg[144][4]  ( .D(\row1_buffer[145][4] ), .CK(clk), .Q(
        \row1_buffer[144][4] ) );
  DFFQXL \row1_buffer_reg[143][4]  ( .D(\row1_buffer[144][4] ), .CK(clk), .Q(
        \row1_buffer[143][4] ) );
  DFFQXL \row1_buffer_reg[142][4]  ( .D(\row1_buffer[143][4] ), .CK(clk), .Q(
        \row1_buffer[142][4] ) );
  DFFQXL \row1_buffer_reg[141][4]  ( .D(\row1_buffer[142][4] ), .CK(clk), .Q(
        \row1_buffer[141][4] ) );
  DFFQXL \row1_buffer_reg[140][4]  ( .D(\row1_buffer[141][4] ), .CK(clk), .Q(
        \row1_buffer[140][4] ) );
  DFFQXL \row1_buffer_reg[139][4]  ( .D(\row1_buffer[140][4] ), .CK(clk), .Q(
        \row1_buffer[139][4] ) );
  DFFQXL \row1_buffer_reg[138][4]  ( .D(\row1_buffer[139][4] ), .CK(clk), .Q(
        \row1_buffer[138][4] ) );
  DFFQXL \row1_buffer_reg[137][4]  ( .D(\row1_buffer[138][4] ), .CK(clk), .Q(
        \row1_buffer[137][4] ) );
  DFFQXL \row1_buffer_reg[136][4]  ( .D(\row1_buffer[137][4] ), .CK(clk), .Q(
        \row1_buffer[136][4] ) );
  DFFQXL \row1_buffer_reg[135][4]  ( .D(\row1_buffer[136][4] ), .CK(clk), .Q(
        \row1_buffer[135][4] ) );
  DFFQXL \row1_buffer_reg[134][4]  ( .D(\row1_buffer[135][4] ), .CK(clk), .Q(
        \row1_buffer[134][4] ) );
  DFFQXL \row1_buffer_reg[133][4]  ( .D(\row1_buffer[134][4] ), .CK(clk), .Q(
        \row1_buffer[133][4] ) );
  DFFQXL \row1_buffer_reg[132][4]  ( .D(\row1_buffer[133][4] ), .CK(clk), .Q(
        \row1_buffer[132][4] ) );
  DFFQXL \row1_buffer_reg[131][4]  ( .D(\row1_buffer[132][4] ), .CK(clk), .Q(
        \row1_buffer[131][4] ) );
  DFFQXL \row1_buffer_reg[130][4]  ( .D(\row1_buffer[131][4] ), .CK(clk), .Q(
        \row1_buffer[130][4] ) );
  DFFQXL \row1_buffer_reg[129][4]  ( .D(\row1_buffer[130][4] ), .CK(clk), .Q(
        \row1_buffer[129][4] ) );
  DFFQXL \row1_buffer_reg[128][4]  ( .D(\row1_buffer[129][4] ), .CK(clk), .Q(
        \row1_buffer[128][4] ) );
  DFFQXL \row1_buffer_reg[127][4]  ( .D(\row1_buffer[128][4] ), .CK(clk), .Q(
        \row1_buffer[127][4] ) );
  DFFQXL \row1_buffer_reg[126][4]  ( .D(\row1_buffer[127][4] ), .CK(clk), .Q(
        \row1_buffer[126][4] ) );
  DFFQXL \row1_buffer_reg[125][4]  ( .D(\row1_buffer[126][4] ), .CK(clk), .Q(
        \row1_buffer[125][4] ) );
  DFFQXL \row1_buffer_reg[124][4]  ( .D(\row1_buffer[125][4] ), .CK(clk), .Q(
        \row1_buffer[124][4] ) );
  DFFQXL \row1_buffer_reg[123][4]  ( .D(\row1_buffer[124][4] ), .CK(clk), .Q(
        \row1_buffer[123][4] ) );
  DFFQXL \row1_buffer_reg[122][4]  ( .D(\row1_buffer[123][4] ), .CK(clk), .Q(
        \row1_buffer[122][4] ) );
  DFFQXL \row1_buffer_reg[121][4]  ( .D(\row1_buffer[122][4] ), .CK(clk), .Q(
        \row1_buffer[121][4] ) );
  DFFQXL \row1_buffer_reg[120][4]  ( .D(\row1_buffer[121][4] ), .CK(clk), .Q(
        \row1_buffer[120][4] ) );
  DFFQXL \row1_buffer_reg[119][4]  ( .D(\row1_buffer[120][4] ), .CK(clk), .Q(
        \row1_buffer[119][4] ) );
  DFFQXL \row1_buffer_reg[118][4]  ( .D(\row1_buffer[119][4] ), .CK(clk), .Q(
        \row1_buffer[118][4] ) );
  DFFQXL \row1_buffer_reg[117][4]  ( .D(\row1_buffer[118][4] ), .CK(clk), .Q(
        \row1_buffer[117][4] ) );
  DFFQXL \row1_buffer_reg[116][4]  ( .D(\row1_buffer[117][4] ), .CK(clk), .Q(
        \row1_buffer[116][4] ) );
  DFFQXL \row1_buffer_reg[115][4]  ( .D(\row1_buffer[116][4] ), .CK(clk), .Q(
        \row1_buffer[115][4] ) );
  DFFQXL \row1_buffer_reg[114][4]  ( .D(\row1_buffer[115][4] ), .CK(clk), .Q(
        \row1_buffer[114][4] ) );
  DFFQXL \row1_buffer_reg[113][4]  ( .D(\row1_buffer[114][4] ), .CK(clk), .Q(
        \row1_buffer[113][4] ) );
  DFFQXL \row1_buffer_reg[112][4]  ( .D(\row1_buffer[113][4] ), .CK(clk), .Q(
        \row1_buffer[112][4] ) );
  DFFQXL \row1_buffer_reg[111][4]  ( .D(\row1_buffer[112][4] ), .CK(clk), .Q(
        \row1_buffer[111][4] ) );
  DFFQXL \row1_buffer_reg[110][4]  ( .D(\row1_buffer[111][4] ), .CK(clk), .Q(
        \row1_buffer[110][4] ) );
  DFFQXL \row1_buffer_reg[109][4]  ( .D(\row1_buffer[110][4] ), .CK(clk), .Q(
        \row1_buffer[109][4] ) );
  DFFQXL \row1_buffer_reg[108][4]  ( .D(\row1_buffer[109][4] ), .CK(clk), .Q(
        \row1_buffer[108][4] ) );
  DFFQXL \row1_buffer_reg[107][4]  ( .D(\row1_buffer[108][4] ), .CK(clk), .Q(
        \row1_buffer[107][4] ) );
  DFFQXL \row1_buffer_reg[106][4]  ( .D(\row1_buffer[107][4] ), .CK(clk), .Q(
        \row1_buffer[106][4] ) );
  DFFQXL \row1_buffer_reg[105][4]  ( .D(\row1_buffer[106][4] ), .CK(clk), .Q(
        \row1_buffer[105][4] ) );
  DFFQXL \row1_buffer_reg[104][4]  ( .D(\row1_buffer[105][4] ), .CK(clk), .Q(
        \row1_buffer[104][4] ) );
  DFFQXL \row1_buffer_reg[103][4]  ( .D(\row1_buffer[104][4] ), .CK(clk), .Q(
        \row1_buffer[103][4] ) );
  DFFQXL \row1_buffer_reg[102][4]  ( .D(\row1_buffer[103][4] ), .CK(clk), .Q(
        \row1_buffer[102][4] ) );
  DFFQXL \row1_buffer_reg[101][4]  ( .D(\row1_buffer[102][4] ), .CK(clk), .Q(
        \row1_buffer[101][4] ) );
  DFFQXL \row1_buffer_reg[100][4]  ( .D(\row1_buffer[101][4] ), .CK(clk), .Q(
        \row1_buffer[100][4] ) );
  DFFQXL \row1_buffer_reg[99][4]  ( .D(\row1_buffer[100][4] ), .CK(clk), .Q(
        \row1_buffer[99][4] ) );
  DFFQXL \row1_buffer_reg[98][4]  ( .D(\row1_buffer[99][4] ), .CK(clk), .Q(
        \row1_buffer[98][4] ) );
  DFFQXL \row1_buffer_reg[97][4]  ( .D(\row1_buffer[98][4] ), .CK(clk), .Q(
        \row1_buffer[97][4] ) );
  DFFQXL \row1_buffer_reg[96][4]  ( .D(\row1_buffer[97][4] ), .CK(clk), .Q(
        \row1_buffer[96][4] ) );
  DFFQXL \row1_buffer_reg[95][4]  ( .D(\row1_buffer[96][4] ), .CK(clk), .Q(
        \row1_buffer[95][4] ) );
  DFFQXL \row1_buffer_reg[94][4]  ( .D(\row1_buffer[95][4] ), .CK(clk), .Q(
        \row1_buffer[94][4] ) );
  DFFQXL \row1_buffer_reg[93][4]  ( .D(\row1_buffer[94][4] ), .CK(clk), .Q(
        \row1_buffer[93][4] ) );
  DFFQXL \row1_buffer_reg[92][4]  ( .D(\row1_buffer[93][4] ), .CK(clk), .Q(
        \row1_buffer[92][4] ) );
  DFFQXL \row1_buffer_reg[91][4]  ( .D(\row1_buffer[92][4] ), .CK(clk), .Q(
        \row1_buffer[91][4] ) );
  DFFQXL \row1_buffer_reg[90][4]  ( .D(\row1_buffer[91][4] ), .CK(clk), .Q(
        \row1_buffer[90][4] ) );
  DFFQXL \row1_buffer_reg[89][4]  ( .D(\row1_buffer[90][4] ), .CK(clk), .Q(
        \row1_buffer[89][4] ) );
  DFFQXL \row1_buffer_reg[88][4]  ( .D(\row1_buffer[89][4] ), .CK(clk), .Q(
        \row1_buffer[88][4] ) );
  DFFQXL \row1_buffer_reg[87][4]  ( .D(\row1_buffer[88][4] ), .CK(clk), .Q(
        \row1_buffer[87][4] ) );
  DFFQXL \row1_buffer_reg[86][4]  ( .D(\row1_buffer[87][4] ), .CK(clk), .Q(
        \row1_buffer[86][4] ) );
  DFFQXL \row1_buffer_reg[85][4]  ( .D(\row1_buffer[86][4] ), .CK(clk), .Q(
        \row1_buffer[85][4] ) );
  DFFQXL \row1_buffer_reg[84][4]  ( .D(\row1_buffer[85][4] ), .CK(clk), .Q(
        \row1_buffer[84][4] ) );
  DFFQXL \row1_buffer_reg[83][4]  ( .D(\row1_buffer[84][4] ), .CK(clk), .Q(
        \row1_buffer[83][4] ) );
  DFFQXL \row1_buffer_reg[82][4]  ( .D(\row1_buffer[83][4] ), .CK(clk), .Q(
        \row1_buffer[82][4] ) );
  DFFQXL \row1_buffer_reg[81][4]  ( .D(\row1_buffer[82][4] ), .CK(clk), .Q(
        \row1_buffer[81][4] ) );
  DFFQXL \row1_buffer_reg[80][4]  ( .D(\row1_buffer[81][4] ), .CK(clk), .Q(
        \row1_buffer[80][4] ) );
  DFFQXL \row1_buffer_reg[79][4]  ( .D(\row1_buffer[80][4] ), .CK(clk), .Q(
        \row1_buffer[79][4] ) );
  DFFQXL \row1_buffer_reg[78][4]  ( .D(\row1_buffer[79][4] ), .CK(clk), .Q(
        \row1_buffer[78][4] ) );
  DFFQXL \row1_buffer_reg[77][4]  ( .D(\row1_buffer[78][4] ), .CK(clk), .Q(
        \row1_buffer[77][4] ) );
  DFFQXL \row1_buffer_reg[76][4]  ( .D(\row1_buffer[77][4] ), .CK(clk), .Q(
        \row1_buffer[76][4] ) );
  DFFQXL \row1_buffer_reg[75][4]  ( .D(\row1_buffer[76][4] ), .CK(clk), .Q(
        \row1_buffer[75][4] ) );
  DFFQXL \row1_buffer_reg[74][4]  ( .D(\row1_buffer[75][4] ), .CK(clk), .Q(
        \row1_buffer[74][4] ) );
  DFFQXL \row1_buffer_reg[73][4]  ( .D(\row1_buffer[74][4] ), .CK(clk), .Q(
        \row1_buffer[73][4] ) );
  DFFQXL \row1_buffer_reg[72][4]  ( .D(\row1_buffer[73][4] ), .CK(clk), .Q(
        \row1_buffer[72][4] ) );
  DFFQXL \row1_buffer_reg[71][4]  ( .D(\row1_buffer[72][4] ), .CK(clk), .Q(
        \row1_buffer[71][4] ) );
  DFFQXL \row1_buffer_reg[70][4]  ( .D(\row1_buffer[71][4] ), .CK(clk), .Q(
        \row1_buffer[70][4] ) );
  DFFQXL \row1_buffer_reg[69][4]  ( .D(\row1_buffer[70][4] ), .CK(clk), .Q(
        \row1_buffer[69][4] ) );
  DFFQXL \row1_buffer_reg[68][4]  ( .D(\row1_buffer[69][4] ), .CK(clk), .Q(
        \row1_buffer[68][4] ) );
  DFFQXL \row1_buffer_reg[67][4]  ( .D(\row1_buffer[68][4] ), .CK(clk), .Q(
        \row1_buffer[67][4] ) );
  DFFQXL \row1_buffer_reg[66][4]  ( .D(\row1_buffer[67][4] ), .CK(clk), .Q(
        \row1_buffer[66][4] ) );
  DFFQXL \row1_buffer_reg[65][4]  ( .D(\row1_buffer[66][4] ), .CK(clk), .Q(
        \row1_buffer[65][4] ) );
  DFFQXL \row1_buffer_reg[64][4]  ( .D(\row1_buffer[65][4] ), .CK(clk), .Q(
        \row1_buffer[64][4] ) );
  DFFQXL \row1_buffer_reg[63][4]  ( .D(\row1_buffer[64][4] ), .CK(clk), .Q(
        \row1_buffer[63][4] ) );
  DFFQXL \row1_buffer_reg[62][4]  ( .D(\row1_buffer[63][4] ), .CK(clk), .Q(
        \row1_buffer[62][4] ) );
  DFFQXL \row1_buffer_reg[61][4]  ( .D(\row1_buffer[62][4] ), .CK(clk), .Q(
        \row1_buffer[61][4] ) );
  DFFQXL \row1_buffer_reg[60][4]  ( .D(\row1_buffer[61][4] ), .CK(clk), .Q(
        \row1_buffer[60][4] ) );
  DFFQXL \row1_buffer_reg[59][4]  ( .D(\row1_buffer[60][4] ), .CK(clk), .Q(
        \row1_buffer[59][4] ) );
  DFFQXL \row1_buffer_reg[58][4]  ( .D(\row1_buffer[59][4] ), .CK(clk), .Q(
        \row1_buffer[58][4] ) );
  DFFQXL \row1_buffer_reg[57][4]  ( .D(\row1_buffer[58][4] ), .CK(clk), .Q(
        \row1_buffer[57][4] ) );
  DFFQXL \row1_buffer_reg[56][4]  ( .D(\row1_buffer[57][4] ), .CK(clk), .Q(
        \row1_buffer[56][4] ) );
  DFFQXL \row1_buffer_reg[55][4]  ( .D(\row1_buffer[56][4] ), .CK(clk), .Q(
        \row1_buffer[55][4] ) );
  DFFQXL \row1_buffer_reg[54][4]  ( .D(\row1_buffer[55][4] ), .CK(clk), .Q(
        \row1_buffer[54][4] ) );
  DFFQXL \row1_buffer_reg[53][4]  ( .D(\row1_buffer[54][4] ), .CK(clk), .Q(
        \row1_buffer[53][4] ) );
  DFFQXL \row1_buffer_reg[52][4]  ( .D(\row1_buffer[53][4] ), .CK(clk), .Q(
        \row1_buffer[52][4] ) );
  DFFQXL \row1_buffer_reg[51][4]  ( .D(\row1_buffer[52][4] ), .CK(clk), .Q(
        \row1_buffer[51][4] ) );
  DFFQXL \row1_buffer_reg[50][4]  ( .D(\row1_buffer[51][4] ), .CK(clk), .Q(
        \row1_buffer[50][4] ) );
  DFFQXL \row1_buffer_reg[49][4]  ( .D(\row1_buffer[50][4] ), .CK(clk), .Q(
        \row1_buffer[49][4] ) );
  DFFQXL \row1_buffer_reg[48][4]  ( .D(\row1_buffer[49][4] ), .CK(clk), .Q(
        \row1_buffer[48][4] ) );
  DFFQXL \row1_buffer_reg[47][4]  ( .D(\row1_buffer[48][4] ), .CK(clk), .Q(
        \row1_buffer[47][4] ) );
  DFFQXL \row1_buffer_reg[46][4]  ( .D(\row1_buffer[47][4] ), .CK(clk), .Q(
        \row1_buffer[46][4] ) );
  DFFQXL \row1_buffer_reg[45][4]  ( .D(\row1_buffer[46][4] ), .CK(clk), .Q(
        \row1_buffer[45][4] ) );
  DFFQXL \row1_buffer_reg[44][4]  ( .D(\row1_buffer[45][4] ), .CK(clk), .Q(
        \row1_buffer[44][4] ) );
  DFFQXL \row1_buffer_reg[43][4]  ( .D(\row1_buffer[44][4] ), .CK(clk), .Q(
        \row1_buffer[43][4] ) );
  DFFQXL \row1_buffer_reg[42][4]  ( .D(\row1_buffer[43][4] ), .CK(clk), .Q(
        \row1_buffer[42][4] ) );
  DFFQXL \row1_buffer_reg[41][4]  ( .D(\row1_buffer[42][4] ), .CK(clk), .Q(
        \row1_buffer[41][4] ) );
  DFFQXL \row1_buffer_reg[40][4]  ( .D(\row1_buffer[41][4] ), .CK(clk), .Q(
        \row1_buffer[40][4] ) );
  DFFQXL \row1_buffer_reg[39][4]  ( .D(\row1_buffer[40][4] ), .CK(clk), .Q(
        \row1_buffer[39][4] ) );
  DFFQXL \row1_buffer_reg[38][4]  ( .D(\row1_buffer[39][4] ), .CK(clk), .Q(
        \row1_buffer[38][4] ) );
  DFFQXL \row1_buffer_reg[37][4]  ( .D(\row1_buffer[38][4] ), .CK(clk), .Q(
        \row1_buffer[37][4] ) );
  DFFQXL \row1_buffer_reg[36][4]  ( .D(\row1_buffer[37][4] ), .CK(clk), .Q(
        \row1_buffer[36][4] ) );
  DFFQXL \row1_buffer_reg[35][4]  ( .D(\row1_buffer[36][4] ), .CK(clk), .Q(
        \row1_buffer[35][4] ) );
  DFFQXL \row1_buffer_reg[34][4]  ( .D(\row1_buffer[35][4] ), .CK(clk), .Q(
        \row1_buffer[34][4] ) );
  DFFQXL \row1_buffer_reg[33][4]  ( .D(\row1_buffer[34][4] ), .CK(clk), .Q(
        \row1_buffer[33][4] ) );
  DFFQXL \row1_buffer_reg[32][4]  ( .D(\row1_buffer[33][4] ), .CK(clk), .Q(
        \row1_buffer[32][4] ) );
  DFFQXL \row1_buffer_reg[31][4]  ( .D(\row1_buffer[32][4] ), .CK(clk), .Q(
        \row1_buffer[31][4] ) );
  DFFQXL \row1_buffer_reg[30][4]  ( .D(\row1_buffer[31][4] ), .CK(clk), .Q(
        \row1_buffer[30][4] ) );
  DFFQXL \row1_buffer_reg[29][4]  ( .D(\row1_buffer[30][4] ), .CK(clk), .Q(
        \row1_buffer[29][4] ) );
  DFFQXL \row1_buffer_reg[28][4]  ( .D(\row1_buffer[29][4] ), .CK(clk), .Q(
        \row1_buffer[28][4] ) );
  DFFQXL \row1_buffer_reg[27][4]  ( .D(\row1_buffer[28][4] ), .CK(clk), .Q(
        \row1_buffer[27][4] ) );
  DFFQXL \row1_buffer_reg[26][4]  ( .D(\row1_buffer[27][4] ), .CK(clk), .Q(
        \row1_buffer[26][4] ) );
  DFFQXL \row1_buffer_reg[25][4]  ( .D(\row1_buffer[26][4] ), .CK(clk), .Q(
        \row1_buffer[25][4] ) );
  DFFQXL \row1_buffer_reg[24][4]  ( .D(\row1_buffer[25][4] ), .CK(clk), .Q(
        \row1_buffer[24][4] ) );
  DFFQXL \row1_buffer_reg[23][4]  ( .D(\row1_buffer[24][4] ), .CK(clk), .Q(
        \row1_buffer[23][4] ) );
  DFFQXL \row1_buffer_reg[22][4]  ( .D(\row1_buffer[23][4] ), .CK(clk), .Q(
        \row1_buffer[22][4] ) );
  DFFQXL \row1_buffer_reg[21][4]  ( .D(\row1_buffer[22][4] ), .CK(clk), .Q(
        \row1_buffer[21][4] ) );
  DFFQXL \row1_buffer_reg[20][4]  ( .D(\row1_buffer[21][4] ), .CK(clk), .Q(
        \row1_buffer[20][4] ) );
  DFFQXL \row1_buffer_reg[19][4]  ( .D(\row1_buffer[20][4] ), .CK(clk), .Q(
        \row1_buffer[19][4] ) );
  DFFQXL \row1_buffer_reg[18][4]  ( .D(\row1_buffer[19][4] ), .CK(clk), .Q(
        \row1_buffer[18][4] ) );
  DFFQXL \row1_buffer_reg[17][4]  ( .D(\row1_buffer[18][4] ), .CK(clk), .Q(
        \row1_buffer[17][4] ) );
  DFFQXL \row1_buffer_reg[16][4]  ( .D(\row1_buffer[17][4] ), .CK(clk), .Q(
        \row1_buffer[16][4] ) );
  DFFQXL \row1_buffer_reg[15][4]  ( .D(\row1_buffer[16][4] ), .CK(clk), .Q(
        \row1_buffer[15][4] ) );
  DFFQXL \row1_buffer_reg[14][4]  ( .D(\row1_buffer[15][4] ), .CK(clk), .Q(
        \row1_buffer[14][4] ) );
  DFFQXL \row1_buffer_reg[13][4]  ( .D(\row1_buffer[14][4] ), .CK(clk), .Q(
        \row1_buffer[13][4] ) );
  DFFQXL \row1_buffer_reg[12][4]  ( .D(\row1_buffer[13][4] ), .CK(clk), .Q(
        \row1_buffer[12][4] ) );
  DFFQXL \row1_buffer_reg[11][4]  ( .D(\row1_buffer[12][4] ), .CK(clk), .Q(
        \row1_buffer[11][4] ) );
  DFFQXL \row1_buffer_reg[10][4]  ( .D(\row1_buffer[11][4] ), .CK(clk), .Q(
        \row1_buffer[10][4] ) );
  DFFQXL \row1_buffer_reg[9][4]  ( .D(\row1_buffer[10][4] ), .CK(clk), .Q(
        \row1_buffer[9][4] ) );
  DFFQXL \row1_buffer_reg[8][4]  ( .D(\row1_buffer[9][4] ), .CK(clk), .Q(
        \row1_buffer[8][4] ) );
  DFFQXL \row1_buffer_reg[7][4]  ( .D(\row1_buffer[8][4] ), .CK(clk), .Q(
        \row1_buffer[7][4] ) );
  DFFQXL \row1_buffer_reg[6][4]  ( .D(\row1_buffer[7][4] ), .CK(clk), .Q(
        \row1_buffer[6][4] ) );
  DFFQXL \row1_buffer_reg[5][4]  ( .D(\row1_buffer[6][4] ), .CK(clk), .Q(
        \row1_buffer[5][4] ) );
  DFFQXL \row1_buffer_reg[4][4]  ( .D(\row1_buffer[5][4] ), .CK(clk), .Q(
        \row1_buffer[4][4] ) );
  DFFQXL \row1_buffer_reg[3][4]  ( .D(\row1_buffer[4][4] ), .CK(clk), .Q(
        \row1_buffer[3][4] ) );
  DFFQXL \row2_buffer_reg[225][3]  ( .D(\row3_buffer[0][3] ), .CK(clk), .Q(
        \row2_buffer[225][3] ) );
  DFFQXL \row2_buffer_reg[224][3]  ( .D(\row2_buffer[225][3] ), .CK(clk), .Q(
        \row2_buffer[224][3] ) );
  DFFQXL \row2_buffer_reg[223][3]  ( .D(\row2_buffer[224][3] ), .CK(clk), .Q(
        \row2_buffer[223][3] ) );
  DFFQXL \row2_buffer_reg[222][3]  ( .D(\row2_buffer[223][3] ), .CK(clk), .Q(
        \row2_buffer[222][3] ) );
  DFFQXL \row2_buffer_reg[221][3]  ( .D(\row2_buffer[222][3] ), .CK(clk), .Q(
        \row2_buffer[221][3] ) );
  DFFQXL \row2_buffer_reg[220][3]  ( .D(\row2_buffer[221][3] ), .CK(clk), .Q(
        \row2_buffer[220][3] ) );
  DFFQXL \row2_buffer_reg[219][3]  ( .D(\row2_buffer[220][3] ), .CK(clk), .Q(
        \row2_buffer[219][3] ) );
  DFFQXL \row2_buffer_reg[218][3]  ( .D(\row2_buffer[219][3] ), .CK(clk), .Q(
        \row2_buffer[218][3] ) );
  DFFQXL \row2_buffer_reg[217][3]  ( .D(\row2_buffer[218][3] ), .CK(clk), .Q(
        \row2_buffer[217][3] ) );
  DFFQXL \row2_buffer_reg[216][3]  ( .D(\row2_buffer[217][3] ), .CK(clk), .Q(
        \row2_buffer[216][3] ) );
  DFFQXL \row2_buffer_reg[215][3]  ( .D(\row2_buffer[216][3] ), .CK(clk), .Q(
        \row2_buffer[215][3] ) );
  DFFQXL \row2_buffer_reg[214][3]  ( .D(\row2_buffer[215][3] ), .CK(clk), .Q(
        \row2_buffer[214][3] ) );
  DFFQXL \row2_buffer_reg[213][3]  ( .D(\row2_buffer[214][3] ), .CK(clk), .Q(
        \row2_buffer[213][3] ) );
  DFFQXL \row2_buffer_reg[212][3]  ( .D(\row2_buffer[213][3] ), .CK(clk), .Q(
        \row2_buffer[212][3] ) );
  DFFQXL \row2_buffer_reg[211][3]  ( .D(\row2_buffer[212][3] ), .CK(clk), .Q(
        \row2_buffer[211][3] ) );
  DFFQXL \row2_buffer_reg[210][3]  ( .D(\row2_buffer[211][3] ), .CK(clk), .Q(
        \row2_buffer[210][3] ) );
  DFFQXL \row2_buffer_reg[209][3]  ( .D(\row2_buffer[210][3] ), .CK(clk), .Q(
        \row2_buffer[209][3] ) );
  DFFQXL \row2_buffer_reg[208][3]  ( .D(\row2_buffer[209][3] ), .CK(clk), .Q(
        \row2_buffer[208][3] ) );
  DFFQXL \row2_buffer_reg[207][3]  ( .D(\row2_buffer[208][3] ), .CK(clk), .Q(
        \row2_buffer[207][3] ) );
  DFFQXL \row2_buffer_reg[206][3]  ( .D(\row2_buffer[207][3] ), .CK(clk), .Q(
        \row2_buffer[206][3] ) );
  DFFQXL \row2_buffer_reg[205][3]  ( .D(\row2_buffer[206][3] ), .CK(clk), .Q(
        \row2_buffer[205][3] ) );
  DFFQXL \row2_buffer_reg[204][3]  ( .D(\row2_buffer[205][3] ), .CK(clk), .Q(
        \row2_buffer[204][3] ) );
  DFFQXL \row2_buffer_reg[203][3]  ( .D(\row2_buffer[204][3] ), .CK(clk), .Q(
        \row2_buffer[203][3] ) );
  DFFQXL \row2_buffer_reg[202][3]  ( .D(\row2_buffer[203][3] ), .CK(clk), .Q(
        \row2_buffer[202][3] ) );
  DFFQXL \row2_buffer_reg[201][3]  ( .D(\row2_buffer[202][3] ), .CK(clk), .Q(
        \row2_buffer[201][3] ) );
  DFFQXL \row2_buffer_reg[200][3]  ( .D(\row2_buffer[201][3] ), .CK(clk), .Q(
        \row2_buffer[200][3] ) );
  DFFQXL \row2_buffer_reg[199][3]  ( .D(\row2_buffer[200][3] ), .CK(clk), .Q(
        \row2_buffer[199][3] ) );
  DFFQXL \row2_buffer_reg[198][3]  ( .D(\row2_buffer[199][3] ), .CK(clk), .Q(
        \row2_buffer[198][3] ) );
  DFFQXL \row2_buffer_reg[197][3]  ( .D(\row2_buffer[198][3] ), .CK(clk), .Q(
        \row2_buffer[197][3] ) );
  DFFQXL \row2_buffer_reg[196][3]  ( .D(\row2_buffer[197][3] ), .CK(clk), .Q(
        \row2_buffer[196][3] ) );
  DFFQXL \row2_buffer_reg[195][3]  ( .D(\row2_buffer[196][3] ), .CK(clk), .Q(
        \row2_buffer[195][3] ) );
  DFFQXL \row2_buffer_reg[194][3]  ( .D(\row2_buffer[195][3] ), .CK(clk), .Q(
        \row2_buffer[194][3] ) );
  DFFQXL \row2_buffer_reg[193][3]  ( .D(\row2_buffer[194][3] ), .CK(clk), .Q(
        \row2_buffer[193][3] ) );
  DFFQXL \row2_buffer_reg[192][3]  ( .D(\row2_buffer[193][3] ), .CK(clk), .Q(
        \row2_buffer[192][3] ) );
  DFFQXL \row2_buffer_reg[191][3]  ( .D(\row2_buffer[192][3] ), .CK(clk), .Q(
        \row2_buffer[191][3] ) );
  DFFQXL \row2_buffer_reg[190][3]  ( .D(\row2_buffer[191][3] ), .CK(clk), .Q(
        \row2_buffer[190][3] ) );
  DFFQXL \row2_buffer_reg[189][3]  ( .D(\row2_buffer[190][3] ), .CK(clk), .Q(
        \row2_buffer[189][3] ) );
  DFFQXL \row2_buffer_reg[188][3]  ( .D(\row2_buffer[189][3] ), .CK(clk), .Q(
        \row2_buffer[188][3] ) );
  DFFQXL \row2_buffer_reg[187][3]  ( .D(\row2_buffer[188][3] ), .CK(clk), .Q(
        \row2_buffer[187][3] ) );
  DFFQXL \row2_buffer_reg[186][3]  ( .D(\row2_buffer[187][3] ), .CK(clk), .Q(
        \row2_buffer[186][3] ) );
  DFFQXL \row2_buffer_reg[185][3]  ( .D(\row2_buffer[186][3] ), .CK(clk), .Q(
        \row2_buffer[185][3] ) );
  DFFQXL \row2_buffer_reg[184][3]  ( .D(\row2_buffer[185][3] ), .CK(clk), .Q(
        \row2_buffer[184][3] ) );
  DFFQXL \row2_buffer_reg[183][3]  ( .D(\row2_buffer[184][3] ), .CK(clk), .Q(
        \row2_buffer[183][3] ) );
  DFFQXL \row2_buffer_reg[182][3]  ( .D(\row2_buffer[183][3] ), .CK(clk), .Q(
        \row2_buffer[182][3] ) );
  DFFQXL \row2_buffer_reg[181][3]  ( .D(\row2_buffer[182][3] ), .CK(clk), .Q(
        \row2_buffer[181][3] ) );
  DFFQXL \row2_buffer_reg[180][3]  ( .D(\row2_buffer[181][3] ), .CK(clk), .Q(
        \row2_buffer[180][3] ) );
  DFFQXL \row2_buffer_reg[179][3]  ( .D(\row2_buffer[180][3] ), .CK(clk), .Q(
        \row2_buffer[179][3] ) );
  DFFQXL \row2_buffer_reg[178][3]  ( .D(\row2_buffer[179][3] ), .CK(clk), .Q(
        \row2_buffer[178][3] ) );
  DFFQXL \row2_buffer_reg[177][3]  ( .D(\row2_buffer[178][3] ), .CK(clk), .Q(
        \row2_buffer[177][3] ) );
  DFFQXL \row2_buffer_reg[176][3]  ( .D(\row2_buffer[177][3] ), .CK(clk), .Q(
        \row2_buffer[176][3] ) );
  DFFQXL \row2_buffer_reg[175][3]  ( .D(\row2_buffer[176][3] ), .CK(clk), .Q(
        \row2_buffer[175][3] ) );
  DFFQXL \row2_buffer_reg[174][3]  ( .D(\row2_buffer[175][3] ), .CK(clk), .Q(
        \row2_buffer[174][3] ) );
  DFFQXL \row2_buffer_reg[173][3]  ( .D(\row2_buffer[174][3] ), .CK(clk), .Q(
        \row2_buffer[173][3] ) );
  DFFQXL \row2_buffer_reg[172][3]  ( .D(\row2_buffer[173][3] ), .CK(clk), .Q(
        \row2_buffer[172][3] ) );
  DFFQXL \row2_buffer_reg[171][3]  ( .D(\row2_buffer[172][3] ), .CK(clk), .Q(
        \row2_buffer[171][3] ) );
  DFFQXL \row2_buffer_reg[170][3]  ( .D(\row2_buffer[171][3] ), .CK(clk), .Q(
        \row2_buffer[170][3] ) );
  DFFQXL \row2_buffer_reg[169][3]  ( .D(\row2_buffer[170][3] ), .CK(clk), .Q(
        \row2_buffer[169][3] ) );
  DFFQXL \row2_buffer_reg[168][3]  ( .D(\row2_buffer[169][3] ), .CK(clk), .Q(
        \row2_buffer[168][3] ) );
  DFFQXL \row2_buffer_reg[167][3]  ( .D(\row2_buffer[168][3] ), .CK(clk), .Q(
        \row2_buffer[167][3] ) );
  DFFQXL \row2_buffer_reg[166][3]  ( .D(\row2_buffer[167][3] ), .CK(clk), .Q(
        \row2_buffer[166][3] ) );
  DFFQXL \row2_buffer_reg[165][3]  ( .D(\row2_buffer[166][3] ), .CK(clk), .Q(
        \row2_buffer[165][3] ) );
  DFFQXL \row2_buffer_reg[164][3]  ( .D(\row2_buffer[165][3] ), .CK(clk), .Q(
        \row2_buffer[164][3] ) );
  DFFQXL \row2_buffer_reg[163][3]  ( .D(\row2_buffer[164][3] ), .CK(clk), .Q(
        \row2_buffer[163][3] ) );
  DFFQXL \row2_buffer_reg[162][3]  ( .D(\row2_buffer[163][3] ), .CK(clk), .Q(
        \row2_buffer[162][3] ) );
  DFFQXL \row2_buffer_reg[161][3]  ( .D(\row2_buffer[162][3] ), .CK(clk), .Q(
        \row2_buffer[161][3] ) );
  DFFQXL \row2_buffer_reg[160][3]  ( .D(\row2_buffer[161][3] ), .CK(clk), .Q(
        \row2_buffer[160][3] ) );
  DFFQXL \row2_buffer_reg[159][3]  ( .D(\row2_buffer[160][3] ), .CK(clk), .Q(
        \row2_buffer[159][3] ) );
  DFFQXL \row2_buffer_reg[158][3]  ( .D(\row2_buffer[159][3] ), .CK(clk), .Q(
        \row2_buffer[158][3] ) );
  DFFQXL \row2_buffer_reg[157][3]  ( .D(\row2_buffer[158][3] ), .CK(clk), .Q(
        \row2_buffer[157][3] ) );
  DFFQXL \row2_buffer_reg[156][3]  ( .D(\row2_buffer[157][3] ), .CK(clk), .Q(
        \row2_buffer[156][3] ) );
  DFFQXL \row2_buffer_reg[155][3]  ( .D(\row2_buffer[156][3] ), .CK(clk), .Q(
        \row2_buffer[155][3] ) );
  DFFQXL \row2_buffer_reg[154][3]  ( .D(\row2_buffer[155][3] ), .CK(clk), .Q(
        \row2_buffer[154][3] ) );
  DFFQXL \row2_buffer_reg[153][3]  ( .D(\row2_buffer[154][3] ), .CK(clk), .Q(
        \row2_buffer[153][3] ) );
  DFFQXL \row2_buffer_reg[152][3]  ( .D(\row2_buffer[153][3] ), .CK(clk), .Q(
        \row2_buffer[152][3] ) );
  DFFQXL \row2_buffer_reg[151][3]  ( .D(\row2_buffer[152][3] ), .CK(clk), .Q(
        \row2_buffer[151][3] ) );
  DFFQXL \row2_buffer_reg[150][3]  ( .D(\row2_buffer[151][3] ), .CK(clk), .Q(
        \row2_buffer[150][3] ) );
  DFFQXL \row2_buffer_reg[149][3]  ( .D(\row2_buffer[150][3] ), .CK(clk), .Q(
        \row2_buffer[149][3] ) );
  DFFQXL \row2_buffer_reg[148][3]  ( .D(\row2_buffer[149][3] ), .CK(clk), .Q(
        \row2_buffer[148][3] ) );
  DFFQXL \row2_buffer_reg[147][3]  ( .D(\row2_buffer[148][3] ), .CK(clk), .Q(
        \row2_buffer[147][3] ) );
  DFFQXL \row2_buffer_reg[146][3]  ( .D(\row2_buffer[147][3] ), .CK(clk), .Q(
        \row2_buffer[146][3] ) );
  DFFQXL \row2_buffer_reg[145][3]  ( .D(\row2_buffer[146][3] ), .CK(clk), .Q(
        \row2_buffer[145][3] ) );
  DFFQXL \row2_buffer_reg[144][3]  ( .D(\row2_buffer[145][3] ), .CK(clk), .Q(
        \row2_buffer[144][3] ) );
  DFFQXL \row2_buffer_reg[143][3]  ( .D(\row2_buffer[144][3] ), .CK(clk), .Q(
        \row2_buffer[143][3] ) );
  DFFQXL \row2_buffer_reg[142][3]  ( .D(\row2_buffer[143][3] ), .CK(clk), .Q(
        \row2_buffer[142][3] ) );
  DFFQXL \row2_buffer_reg[141][3]  ( .D(\row2_buffer[142][3] ), .CK(clk), .Q(
        \row2_buffer[141][3] ) );
  DFFQXL \row2_buffer_reg[140][3]  ( .D(\row2_buffer[141][3] ), .CK(clk), .Q(
        \row2_buffer[140][3] ) );
  DFFQXL \row2_buffer_reg[139][3]  ( .D(\row2_buffer[140][3] ), .CK(clk), .Q(
        \row2_buffer[139][3] ) );
  DFFQXL \row2_buffer_reg[138][3]  ( .D(\row2_buffer[139][3] ), .CK(clk), .Q(
        \row2_buffer[138][3] ) );
  DFFQXL \row2_buffer_reg[137][3]  ( .D(\row2_buffer[138][3] ), .CK(clk), .Q(
        \row2_buffer[137][3] ) );
  DFFQXL \row2_buffer_reg[136][3]  ( .D(\row2_buffer[137][3] ), .CK(clk), .Q(
        \row2_buffer[136][3] ) );
  DFFQXL \row2_buffer_reg[135][3]  ( .D(\row2_buffer[136][3] ), .CK(clk), .Q(
        \row2_buffer[135][3] ) );
  DFFQXL \row2_buffer_reg[134][3]  ( .D(\row2_buffer[135][3] ), .CK(clk), .Q(
        \row2_buffer[134][3] ) );
  DFFQXL \row2_buffer_reg[133][3]  ( .D(\row2_buffer[134][3] ), .CK(clk), .Q(
        \row2_buffer[133][3] ) );
  DFFQXL \row2_buffer_reg[132][3]  ( .D(\row2_buffer[133][3] ), .CK(clk), .Q(
        \row2_buffer[132][3] ) );
  DFFQXL \row2_buffer_reg[131][3]  ( .D(\row2_buffer[132][3] ), .CK(clk), .Q(
        \row2_buffer[131][3] ) );
  DFFQXL \row2_buffer_reg[130][3]  ( .D(\row2_buffer[131][3] ), .CK(clk), .Q(
        \row2_buffer[130][3] ) );
  DFFQXL \row2_buffer_reg[129][3]  ( .D(\row2_buffer[130][3] ), .CK(clk), .Q(
        \row2_buffer[129][3] ) );
  DFFQXL \row2_buffer_reg[128][3]  ( .D(\row2_buffer[129][3] ), .CK(clk), .Q(
        \row2_buffer[128][3] ) );
  DFFQXL \row2_buffer_reg[127][3]  ( .D(\row2_buffer[128][3] ), .CK(clk), .Q(
        \row2_buffer[127][3] ) );
  DFFQXL \row2_buffer_reg[126][3]  ( .D(\row2_buffer[127][3] ), .CK(clk), .Q(
        \row2_buffer[126][3] ) );
  DFFQXL \row2_buffer_reg[125][3]  ( .D(\row2_buffer[126][3] ), .CK(clk), .Q(
        \row2_buffer[125][3] ) );
  DFFQXL \row2_buffer_reg[124][3]  ( .D(\row2_buffer[125][3] ), .CK(clk), .Q(
        \row2_buffer[124][3] ) );
  DFFQXL \row2_buffer_reg[123][3]  ( .D(\row2_buffer[124][3] ), .CK(clk), .Q(
        \row2_buffer[123][3] ) );
  DFFQXL \row2_buffer_reg[122][3]  ( .D(\row2_buffer[123][3] ), .CK(clk), .Q(
        \row2_buffer[122][3] ) );
  DFFQXL \row2_buffer_reg[121][3]  ( .D(\row2_buffer[122][3] ), .CK(clk), .Q(
        \row2_buffer[121][3] ) );
  DFFQXL \row2_buffer_reg[120][3]  ( .D(\row2_buffer[121][3] ), .CK(clk), .Q(
        \row2_buffer[120][3] ) );
  DFFQXL \row2_buffer_reg[119][3]  ( .D(\row2_buffer[120][3] ), .CK(clk), .Q(
        \row2_buffer[119][3] ) );
  DFFQXL \row2_buffer_reg[118][3]  ( .D(\row2_buffer[119][3] ), .CK(clk), .Q(
        \row2_buffer[118][3] ) );
  DFFQXL \row2_buffer_reg[117][3]  ( .D(\row2_buffer[118][3] ), .CK(clk), .Q(
        \row2_buffer[117][3] ) );
  DFFQXL \row2_buffer_reg[116][3]  ( .D(\row2_buffer[117][3] ), .CK(clk), .Q(
        \row2_buffer[116][3] ) );
  DFFQXL \row2_buffer_reg[115][3]  ( .D(\row2_buffer[116][3] ), .CK(clk), .Q(
        \row2_buffer[115][3] ) );
  DFFQXL \row2_buffer_reg[114][3]  ( .D(\row2_buffer[115][3] ), .CK(clk), .Q(
        \row2_buffer[114][3] ) );
  DFFQXL \row2_buffer_reg[113][3]  ( .D(\row2_buffer[114][3] ), .CK(clk), .Q(
        \row2_buffer[113][3] ) );
  DFFQXL \row2_buffer_reg[112][3]  ( .D(\row2_buffer[113][3] ), .CK(clk), .Q(
        \row2_buffer[112][3] ) );
  DFFQXL \row2_buffer_reg[111][3]  ( .D(\row2_buffer[112][3] ), .CK(clk), .Q(
        \row2_buffer[111][3] ) );
  DFFQXL \row2_buffer_reg[110][3]  ( .D(\row2_buffer[111][3] ), .CK(clk), .Q(
        \row2_buffer[110][3] ) );
  DFFQXL \row2_buffer_reg[109][3]  ( .D(\row2_buffer[110][3] ), .CK(clk), .Q(
        \row2_buffer[109][3] ) );
  DFFQXL \row2_buffer_reg[108][3]  ( .D(\row2_buffer[109][3] ), .CK(clk), .Q(
        \row2_buffer[108][3] ) );
  DFFQXL \row2_buffer_reg[107][3]  ( .D(\row2_buffer[108][3] ), .CK(clk), .Q(
        \row2_buffer[107][3] ) );
  DFFQXL \row2_buffer_reg[106][3]  ( .D(\row2_buffer[107][3] ), .CK(clk), .Q(
        \row2_buffer[106][3] ) );
  DFFQXL \row2_buffer_reg[105][3]  ( .D(\row2_buffer[106][3] ), .CK(clk), .Q(
        \row2_buffer[105][3] ) );
  DFFQXL \row2_buffer_reg[104][3]  ( .D(\row2_buffer[105][3] ), .CK(clk), .Q(
        \row2_buffer[104][3] ) );
  DFFQXL \row2_buffer_reg[103][3]  ( .D(\row2_buffer[104][3] ), .CK(clk), .Q(
        \row2_buffer[103][3] ) );
  DFFQXL \row2_buffer_reg[102][3]  ( .D(\row2_buffer[103][3] ), .CK(clk), .Q(
        \row2_buffer[102][3] ) );
  DFFQXL \row2_buffer_reg[101][3]  ( .D(\row2_buffer[102][3] ), .CK(clk), .Q(
        \row2_buffer[101][3] ) );
  DFFQXL \row2_buffer_reg[100][3]  ( .D(\row2_buffer[101][3] ), .CK(clk), .Q(
        \row2_buffer[100][3] ) );
  DFFQXL \row2_buffer_reg[99][3]  ( .D(\row2_buffer[100][3] ), .CK(clk), .Q(
        \row2_buffer[99][3] ) );
  DFFQXL \row2_buffer_reg[98][3]  ( .D(\row2_buffer[99][3] ), .CK(clk), .Q(
        \row2_buffer[98][3] ) );
  DFFQXL \row2_buffer_reg[97][3]  ( .D(\row2_buffer[98][3] ), .CK(clk), .Q(
        \row2_buffer[97][3] ) );
  DFFQXL \row2_buffer_reg[96][3]  ( .D(\row2_buffer[97][3] ), .CK(clk), .Q(
        \row2_buffer[96][3] ) );
  DFFQXL \row2_buffer_reg[95][3]  ( .D(\row2_buffer[96][3] ), .CK(clk), .Q(
        \row2_buffer[95][3] ) );
  DFFQXL \row2_buffer_reg[94][3]  ( .D(\row2_buffer[95][3] ), .CK(clk), .Q(
        \row2_buffer[94][3] ) );
  DFFQXL \row2_buffer_reg[93][3]  ( .D(\row2_buffer[94][3] ), .CK(clk), .Q(
        \row2_buffer[93][3] ) );
  DFFQXL \row2_buffer_reg[92][3]  ( .D(\row2_buffer[93][3] ), .CK(clk), .Q(
        \row2_buffer[92][3] ) );
  DFFQXL \row2_buffer_reg[91][3]  ( .D(\row2_buffer[92][3] ), .CK(clk), .Q(
        \row2_buffer[91][3] ) );
  DFFQXL \row2_buffer_reg[90][3]  ( .D(\row2_buffer[91][3] ), .CK(clk), .Q(
        \row2_buffer[90][3] ) );
  DFFQXL \row2_buffer_reg[89][3]  ( .D(\row2_buffer[90][3] ), .CK(clk), .Q(
        \row2_buffer[89][3] ) );
  DFFQXL \row2_buffer_reg[88][3]  ( .D(\row2_buffer[89][3] ), .CK(clk), .Q(
        \row2_buffer[88][3] ) );
  DFFQXL \row2_buffer_reg[87][3]  ( .D(\row2_buffer[88][3] ), .CK(clk), .Q(
        \row2_buffer[87][3] ) );
  DFFQXL \row2_buffer_reg[86][3]  ( .D(\row2_buffer[87][3] ), .CK(clk), .Q(
        \row2_buffer[86][3] ) );
  DFFQXL \row2_buffer_reg[85][3]  ( .D(\row2_buffer[86][3] ), .CK(clk), .Q(
        \row2_buffer[85][3] ) );
  DFFQXL \row2_buffer_reg[84][3]  ( .D(\row2_buffer[85][3] ), .CK(clk), .Q(
        \row2_buffer[84][3] ) );
  DFFQXL \row2_buffer_reg[83][3]  ( .D(\row2_buffer[84][3] ), .CK(clk), .Q(
        \row2_buffer[83][3] ) );
  DFFQXL \row2_buffer_reg[82][3]  ( .D(\row2_buffer[83][3] ), .CK(clk), .Q(
        \row2_buffer[82][3] ) );
  DFFQXL \row2_buffer_reg[81][3]  ( .D(\row2_buffer[82][3] ), .CK(clk), .Q(
        \row2_buffer[81][3] ) );
  DFFQXL \row2_buffer_reg[80][3]  ( .D(\row2_buffer[81][3] ), .CK(clk), .Q(
        \row2_buffer[80][3] ) );
  DFFQXL \row2_buffer_reg[79][3]  ( .D(\row2_buffer[80][3] ), .CK(clk), .Q(
        \row2_buffer[79][3] ) );
  DFFQXL \row2_buffer_reg[78][3]  ( .D(\row2_buffer[79][3] ), .CK(clk), .Q(
        \row2_buffer[78][3] ) );
  DFFQXL \row2_buffer_reg[77][3]  ( .D(\row2_buffer[78][3] ), .CK(clk), .Q(
        \row2_buffer[77][3] ) );
  DFFQXL \row2_buffer_reg[76][3]  ( .D(\row2_buffer[77][3] ), .CK(clk), .Q(
        \row2_buffer[76][3] ) );
  DFFQXL \row2_buffer_reg[75][3]  ( .D(\row2_buffer[76][3] ), .CK(clk), .Q(
        \row2_buffer[75][3] ) );
  DFFQXL \row2_buffer_reg[74][3]  ( .D(\row2_buffer[75][3] ), .CK(clk), .Q(
        \row2_buffer[74][3] ) );
  DFFQXL \row2_buffer_reg[73][3]  ( .D(\row2_buffer[74][3] ), .CK(clk), .Q(
        \row2_buffer[73][3] ) );
  DFFQXL \row2_buffer_reg[72][3]  ( .D(\row2_buffer[73][3] ), .CK(clk), .Q(
        \row2_buffer[72][3] ) );
  DFFQXL \row2_buffer_reg[71][3]  ( .D(\row2_buffer[72][3] ), .CK(clk), .Q(
        \row2_buffer[71][3] ) );
  DFFQXL \row2_buffer_reg[70][3]  ( .D(\row2_buffer[71][3] ), .CK(clk), .Q(
        \row2_buffer[70][3] ) );
  DFFQXL \row2_buffer_reg[69][3]  ( .D(\row2_buffer[70][3] ), .CK(clk), .Q(
        \row2_buffer[69][3] ) );
  DFFQXL \row2_buffer_reg[68][3]  ( .D(\row2_buffer[69][3] ), .CK(clk), .Q(
        \row2_buffer[68][3] ) );
  DFFQXL \row2_buffer_reg[67][3]  ( .D(\row2_buffer[68][3] ), .CK(clk), .Q(
        \row2_buffer[67][3] ) );
  DFFQXL \row2_buffer_reg[66][3]  ( .D(\row2_buffer[67][3] ), .CK(clk), .Q(
        \row2_buffer[66][3] ) );
  DFFQXL \row2_buffer_reg[65][3]  ( .D(\row2_buffer[66][3] ), .CK(clk), .Q(
        \row2_buffer[65][3] ) );
  DFFQXL \row2_buffer_reg[64][3]  ( .D(\row2_buffer[65][3] ), .CK(clk), .Q(
        \row2_buffer[64][3] ) );
  DFFQXL \row2_buffer_reg[63][3]  ( .D(\row2_buffer[64][3] ), .CK(clk), .Q(
        \row2_buffer[63][3] ) );
  DFFQXL \row2_buffer_reg[62][3]  ( .D(\row2_buffer[63][3] ), .CK(clk), .Q(
        \row2_buffer[62][3] ) );
  DFFQXL \row2_buffer_reg[61][3]  ( .D(\row2_buffer[62][3] ), .CK(clk), .Q(
        \row2_buffer[61][3] ) );
  DFFQXL \row2_buffer_reg[60][3]  ( .D(\row2_buffer[61][3] ), .CK(clk), .Q(
        \row2_buffer[60][3] ) );
  DFFQXL \row2_buffer_reg[59][3]  ( .D(\row2_buffer[60][3] ), .CK(clk), .Q(
        \row2_buffer[59][3] ) );
  DFFQXL \row2_buffer_reg[58][3]  ( .D(\row2_buffer[59][3] ), .CK(clk), .Q(
        \row2_buffer[58][3] ) );
  DFFQXL \row2_buffer_reg[57][3]  ( .D(\row2_buffer[58][3] ), .CK(clk), .Q(
        \row2_buffer[57][3] ) );
  DFFQXL \row2_buffer_reg[56][3]  ( .D(\row2_buffer[57][3] ), .CK(clk), .Q(
        \row2_buffer[56][3] ) );
  DFFQXL \row2_buffer_reg[55][3]  ( .D(\row2_buffer[56][3] ), .CK(clk), .Q(
        \row2_buffer[55][3] ) );
  DFFQXL \row2_buffer_reg[54][3]  ( .D(\row2_buffer[55][3] ), .CK(clk), .Q(
        \row2_buffer[54][3] ) );
  DFFQXL \row2_buffer_reg[53][3]  ( .D(\row2_buffer[54][3] ), .CK(clk), .Q(
        \row2_buffer[53][3] ) );
  DFFQXL \row2_buffer_reg[52][3]  ( .D(\row2_buffer[53][3] ), .CK(clk), .Q(
        \row2_buffer[52][3] ) );
  DFFQXL \row2_buffer_reg[51][3]  ( .D(\row2_buffer[52][3] ), .CK(clk), .Q(
        \row2_buffer[51][3] ) );
  DFFQXL \row2_buffer_reg[50][3]  ( .D(\row2_buffer[51][3] ), .CK(clk), .Q(
        \row2_buffer[50][3] ) );
  DFFQXL \row2_buffer_reg[49][3]  ( .D(\row2_buffer[50][3] ), .CK(clk), .Q(
        \row2_buffer[49][3] ) );
  DFFQXL \row2_buffer_reg[48][3]  ( .D(\row2_buffer[49][3] ), .CK(clk), .Q(
        \row2_buffer[48][3] ) );
  DFFQXL \row2_buffer_reg[47][3]  ( .D(\row2_buffer[48][3] ), .CK(clk), .Q(
        \row2_buffer[47][3] ) );
  DFFQXL \row2_buffer_reg[46][3]  ( .D(\row2_buffer[47][3] ), .CK(clk), .Q(
        \row2_buffer[46][3] ) );
  DFFQXL \row2_buffer_reg[45][3]  ( .D(\row2_buffer[46][3] ), .CK(clk), .Q(
        \row2_buffer[45][3] ) );
  DFFQXL \row2_buffer_reg[44][3]  ( .D(\row2_buffer[45][3] ), .CK(clk), .Q(
        \row2_buffer[44][3] ) );
  DFFQXL \row2_buffer_reg[43][3]  ( .D(\row2_buffer[44][3] ), .CK(clk), .Q(
        \row2_buffer[43][3] ) );
  DFFQXL \row2_buffer_reg[42][3]  ( .D(\row2_buffer[43][3] ), .CK(clk), .Q(
        \row2_buffer[42][3] ) );
  DFFQXL \row2_buffer_reg[41][3]  ( .D(\row2_buffer[42][3] ), .CK(clk), .Q(
        \row2_buffer[41][3] ) );
  DFFQXL \row2_buffer_reg[40][3]  ( .D(\row2_buffer[41][3] ), .CK(clk), .Q(
        \row2_buffer[40][3] ) );
  DFFQXL \row2_buffer_reg[39][3]  ( .D(\row2_buffer[40][3] ), .CK(clk), .Q(
        \row2_buffer[39][3] ) );
  DFFQXL \row2_buffer_reg[38][3]  ( .D(\row2_buffer[39][3] ), .CK(clk), .Q(
        \row2_buffer[38][3] ) );
  DFFQXL \row2_buffer_reg[37][3]  ( .D(\row2_buffer[38][3] ), .CK(clk), .Q(
        \row2_buffer[37][3] ) );
  DFFQXL \row2_buffer_reg[36][3]  ( .D(\row2_buffer[37][3] ), .CK(clk), .Q(
        \row2_buffer[36][3] ) );
  DFFQXL \row2_buffer_reg[35][3]  ( .D(\row2_buffer[36][3] ), .CK(clk), .Q(
        \row2_buffer[35][3] ) );
  DFFQXL \row2_buffer_reg[34][3]  ( .D(\row2_buffer[35][3] ), .CK(clk), .Q(
        \row2_buffer[34][3] ) );
  DFFQXL \row2_buffer_reg[33][3]  ( .D(\row2_buffer[34][3] ), .CK(clk), .Q(
        \row2_buffer[33][3] ) );
  DFFQXL \row2_buffer_reg[32][3]  ( .D(\row2_buffer[33][3] ), .CK(clk), .Q(
        \row2_buffer[32][3] ) );
  DFFQXL \row2_buffer_reg[31][3]  ( .D(\row2_buffer[32][3] ), .CK(clk), .Q(
        \row2_buffer[31][3] ) );
  DFFQXL \row2_buffer_reg[30][3]  ( .D(\row2_buffer[31][3] ), .CK(clk), .Q(
        \row2_buffer[30][3] ) );
  DFFQXL \row2_buffer_reg[29][3]  ( .D(\row2_buffer[30][3] ), .CK(clk), .Q(
        \row2_buffer[29][3] ) );
  DFFQXL \row2_buffer_reg[28][3]  ( .D(\row2_buffer[29][3] ), .CK(clk), .Q(
        \row2_buffer[28][3] ) );
  DFFQXL \row2_buffer_reg[27][3]  ( .D(\row2_buffer[28][3] ), .CK(clk), .Q(
        \row2_buffer[27][3] ) );
  DFFQXL \row2_buffer_reg[26][3]  ( .D(\row2_buffer[27][3] ), .CK(clk), .Q(
        \row2_buffer[26][3] ) );
  DFFQXL \row2_buffer_reg[25][3]  ( .D(\row2_buffer[26][3] ), .CK(clk), .Q(
        \row2_buffer[25][3] ) );
  DFFQXL \row2_buffer_reg[24][3]  ( .D(\row2_buffer[25][3] ), .CK(clk), .Q(
        \row2_buffer[24][3] ) );
  DFFQXL \row2_buffer_reg[23][3]  ( .D(\row2_buffer[24][3] ), .CK(clk), .Q(
        \row2_buffer[23][3] ) );
  DFFQXL \row2_buffer_reg[22][3]  ( .D(\row2_buffer[23][3] ), .CK(clk), .Q(
        \row2_buffer[22][3] ) );
  DFFQXL \row2_buffer_reg[21][3]  ( .D(\row2_buffer[22][3] ), .CK(clk), .Q(
        \row2_buffer[21][3] ) );
  DFFQXL \row2_buffer_reg[20][3]  ( .D(\row2_buffer[21][3] ), .CK(clk), .Q(
        \row2_buffer[20][3] ) );
  DFFQXL \row2_buffer_reg[19][3]  ( .D(\row2_buffer[20][3] ), .CK(clk), .Q(
        \row2_buffer[19][3] ) );
  DFFQXL \row2_buffer_reg[18][3]  ( .D(\row2_buffer[19][3] ), .CK(clk), .Q(
        \row2_buffer[18][3] ) );
  DFFQXL \row2_buffer_reg[17][3]  ( .D(\row2_buffer[18][3] ), .CK(clk), .Q(
        \row2_buffer[17][3] ) );
  DFFQXL \row2_buffer_reg[16][3]  ( .D(\row2_buffer[17][3] ), .CK(clk), .Q(
        \row2_buffer[16][3] ) );
  DFFQXL \row2_buffer_reg[15][3]  ( .D(\row2_buffer[16][3] ), .CK(clk), .Q(
        \row2_buffer[15][3] ) );
  DFFQXL \row2_buffer_reg[14][3]  ( .D(\row2_buffer[15][3] ), .CK(clk), .Q(
        \row2_buffer[14][3] ) );
  DFFQXL \row2_buffer_reg[13][3]  ( .D(\row2_buffer[14][3] ), .CK(clk), .Q(
        \row2_buffer[13][3] ) );
  DFFQXL \row2_buffer_reg[12][3]  ( .D(\row2_buffer[13][3] ), .CK(clk), .Q(
        \row2_buffer[12][3] ) );
  DFFQXL \row2_buffer_reg[11][3]  ( .D(\row2_buffer[12][3] ), .CK(clk), .Q(
        \row2_buffer[11][3] ) );
  DFFQXL \row2_buffer_reg[10][3]  ( .D(\row2_buffer[11][3] ), .CK(clk), .Q(
        \row2_buffer[10][3] ) );
  DFFQXL \row2_buffer_reg[9][3]  ( .D(\row2_buffer[10][3] ), .CK(clk), .Q(
        \row2_buffer[9][3] ) );
  DFFQXL \row2_buffer_reg[8][3]  ( .D(\row2_buffer[9][3] ), .CK(clk), .Q(
        \row2_buffer[8][3] ) );
  DFFQXL \row2_buffer_reg[7][3]  ( .D(\row2_buffer[8][3] ), .CK(clk), .Q(
        \row2_buffer[7][3] ) );
  DFFQXL \row2_buffer_reg[6][3]  ( .D(\row2_buffer[7][3] ), .CK(clk), .Q(
        \row2_buffer[6][3] ) );
  DFFQXL \row2_buffer_reg[5][3]  ( .D(\row2_buffer[6][3] ), .CK(clk), .Q(
        \row2_buffer[5][3] ) );
  DFFQXL \row2_buffer_reg[4][3]  ( .D(\row2_buffer[5][3] ), .CK(clk), .Q(
        \row2_buffer[4][3] ) );
  DFFQXL \row2_buffer_reg[3][3]  ( .D(\row2_buffer[4][3] ), .CK(clk), .Q(
        \row2_buffer[3][3] ) );
  DFFQXL \row1_buffer_reg[225][3]  ( .D(\row2_buffer[0][3] ), .CK(clk), .Q(
        \row1_buffer[225][3] ) );
  DFFQXL \row1_buffer_reg[224][3]  ( .D(\row1_buffer[225][3] ), .CK(clk), .Q(
        \row1_buffer[224][3] ) );
  DFFQXL \row1_buffer_reg[223][3]  ( .D(\row1_buffer[224][3] ), .CK(clk), .Q(
        \row1_buffer[223][3] ) );
  DFFQXL \row1_buffer_reg[222][3]  ( .D(\row1_buffer[223][3] ), .CK(clk), .Q(
        \row1_buffer[222][3] ) );
  DFFQXL \row1_buffer_reg[221][3]  ( .D(\row1_buffer[222][3] ), .CK(clk), .Q(
        \row1_buffer[221][3] ) );
  DFFQXL \row1_buffer_reg[220][3]  ( .D(\row1_buffer[221][3] ), .CK(clk), .Q(
        \row1_buffer[220][3] ) );
  DFFQXL \row1_buffer_reg[219][3]  ( .D(\row1_buffer[220][3] ), .CK(clk), .Q(
        \row1_buffer[219][3] ) );
  DFFQXL \row1_buffer_reg[218][3]  ( .D(\row1_buffer[219][3] ), .CK(clk), .Q(
        \row1_buffer[218][3] ) );
  DFFQXL \row1_buffer_reg[217][3]  ( .D(\row1_buffer[218][3] ), .CK(clk), .Q(
        \row1_buffer[217][3] ) );
  DFFQXL \row1_buffer_reg[216][3]  ( .D(\row1_buffer[217][3] ), .CK(clk), .Q(
        \row1_buffer[216][3] ) );
  DFFQXL \row1_buffer_reg[215][3]  ( .D(\row1_buffer[216][3] ), .CK(clk), .Q(
        \row1_buffer[215][3] ) );
  DFFQXL \row1_buffer_reg[214][3]  ( .D(\row1_buffer[215][3] ), .CK(clk), .Q(
        \row1_buffer[214][3] ) );
  DFFQXL \row1_buffer_reg[213][3]  ( .D(\row1_buffer[214][3] ), .CK(clk), .Q(
        \row1_buffer[213][3] ) );
  DFFQXL \row1_buffer_reg[212][3]  ( .D(\row1_buffer[213][3] ), .CK(clk), .Q(
        \row1_buffer[212][3] ) );
  DFFQXL \row1_buffer_reg[211][3]  ( .D(\row1_buffer[212][3] ), .CK(clk), .Q(
        \row1_buffer[211][3] ) );
  DFFQXL \row1_buffer_reg[210][3]  ( .D(\row1_buffer[211][3] ), .CK(clk), .Q(
        \row1_buffer[210][3] ) );
  DFFQXL \row1_buffer_reg[209][3]  ( .D(\row1_buffer[210][3] ), .CK(clk), .Q(
        \row1_buffer[209][3] ) );
  DFFQXL \row1_buffer_reg[208][3]  ( .D(\row1_buffer[209][3] ), .CK(clk), .Q(
        \row1_buffer[208][3] ) );
  DFFQXL \row1_buffer_reg[207][3]  ( .D(\row1_buffer[208][3] ), .CK(clk), .Q(
        \row1_buffer[207][3] ) );
  DFFQXL \row1_buffer_reg[206][3]  ( .D(\row1_buffer[207][3] ), .CK(clk), .Q(
        \row1_buffer[206][3] ) );
  DFFQXL \row1_buffer_reg[205][3]  ( .D(\row1_buffer[206][3] ), .CK(clk), .Q(
        \row1_buffer[205][3] ) );
  DFFQXL \row1_buffer_reg[204][3]  ( .D(\row1_buffer[205][3] ), .CK(clk), .Q(
        \row1_buffer[204][3] ) );
  DFFQXL \row1_buffer_reg[203][3]  ( .D(\row1_buffer[204][3] ), .CK(clk), .Q(
        \row1_buffer[203][3] ) );
  DFFQXL \row1_buffer_reg[202][3]  ( .D(\row1_buffer[203][3] ), .CK(clk), .Q(
        \row1_buffer[202][3] ) );
  DFFQXL \row1_buffer_reg[201][3]  ( .D(\row1_buffer[202][3] ), .CK(clk), .Q(
        \row1_buffer[201][3] ) );
  DFFQXL \row1_buffer_reg[200][3]  ( .D(\row1_buffer[201][3] ), .CK(clk), .Q(
        \row1_buffer[200][3] ) );
  DFFQXL \row1_buffer_reg[199][3]  ( .D(\row1_buffer[200][3] ), .CK(clk), .Q(
        \row1_buffer[199][3] ) );
  DFFQXL \row1_buffer_reg[198][3]  ( .D(\row1_buffer[199][3] ), .CK(clk), .Q(
        \row1_buffer[198][3] ) );
  DFFQXL \row1_buffer_reg[197][3]  ( .D(\row1_buffer[198][3] ), .CK(clk), .Q(
        \row1_buffer[197][3] ) );
  DFFQXL \row1_buffer_reg[196][3]  ( .D(\row1_buffer[197][3] ), .CK(clk), .Q(
        \row1_buffer[196][3] ) );
  DFFQXL \row1_buffer_reg[195][3]  ( .D(\row1_buffer[196][3] ), .CK(clk), .Q(
        \row1_buffer[195][3] ) );
  DFFQXL \row1_buffer_reg[194][3]  ( .D(\row1_buffer[195][3] ), .CK(clk), .Q(
        \row1_buffer[194][3] ) );
  DFFQXL \row1_buffer_reg[193][3]  ( .D(\row1_buffer[194][3] ), .CK(clk), .Q(
        \row1_buffer[193][3] ) );
  DFFQXL \row1_buffer_reg[192][3]  ( .D(\row1_buffer[193][3] ), .CK(clk), .Q(
        \row1_buffer[192][3] ) );
  DFFQXL \row1_buffer_reg[191][3]  ( .D(\row1_buffer[192][3] ), .CK(clk), .Q(
        \row1_buffer[191][3] ) );
  DFFQXL \row1_buffer_reg[190][3]  ( .D(\row1_buffer[191][3] ), .CK(clk), .Q(
        \row1_buffer[190][3] ) );
  DFFQXL \row1_buffer_reg[189][3]  ( .D(\row1_buffer[190][3] ), .CK(clk), .Q(
        \row1_buffer[189][3] ) );
  DFFQXL \row1_buffer_reg[188][3]  ( .D(\row1_buffer[189][3] ), .CK(clk), .Q(
        \row1_buffer[188][3] ) );
  DFFQXL \row1_buffer_reg[187][3]  ( .D(\row1_buffer[188][3] ), .CK(clk), .Q(
        \row1_buffer[187][3] ) );
  DFFQXL \row1_buffer_reg[186][3]  ( .D(\row1_buffer[187][3] ), .CK(clk), .Q(
        \row1_buffer[186][3] ) );
  DFFQXL \row1_buffer_reg[185][3]  ( .D(\row1_buffer[186][3] ), .CK(clk), .Q(
        \row1_buffer[185][3] ) );
  DFFQXL \row1_buffer_reg[184][3]  ( .D(\row1_buffer[185][3] ), .CK(clk), .Q(
        \row1_buffer[184][3] ) );
  DFFQXL \row1_buffer_reg[183][3]  ( .D(\row1_buffer[184][3] ), .CK(clk), .Q(
        \row1_buffer[183][3] ) );
  DFFQXL \row1_buffer_reg[182][3]  ( .D(\row1_buffer[183][3] ), .CK(clk), .Q(
        \row1_buffer[182][3] ) );
  DFFQXL \row1_buffer_reg[181][3]  ( .D(\row1_buffer[182][3] ), .CK(clk), .Q(
        \row1_buffer[181][3] ) );
  DFFQXL \row1_buffer_reg[180][3]  ( .D(\row1_buffer[181][3] ), .CK(clk), .Q(
        \row1_buffer[180][3] ) );
  DFFQXL \row1_buffer_reg[179][3]  ( .D(\row1_buffer[180][3] ), .CK(clk), .Q(
        \row1_buffer[179][3] ) );
  DFFQXL \row1_buffer_reg[178][3]  ( .D(\row1_buffer[179][3] ), .CK(clk), .Q(
        \row1_buffer[178][3] ) );
  DFFQXL \row1_buffer_reg[177][3]  ( .D(\row1_buffer[178][3] ), .CK(clk), .Q(
        \row1_buffer[177][3] ) );
  DFFQXL \row1_buffer_reg[176][3]  ( .D(\row1_buffer[177][3] ), .CK(clk), .Q(
        \row1_buffer[176][3] ) );
  DFFQXL \row1_buffer_reg[175][3]  ( .D(\row1_buffer[176][3] ), .CK(clk), .Q(
        \row1_buffer[175][3] ) );
  DFFQXL \row1_buffer_reg[174][3]  ( .D(\row1_buffer[175][3] ), .CK(clk), .Q(
        \row1_buffer[174][3] ) );
  DFFQXL \row1_buffer_reg[173][3]  ( .D(\row1_buffer[174][3] ), .CK(clk), .Q(
        \row1_buffer[173][3] ) );
  DFFQXL \row1_buffer_reg[172][3]  ( .D(\row1_buffer[173][3] ), .CK(clk), .Q(
        \row1_buffer[172][3] ) );
  DFFQXL \row1_buffer_reg[171][3]  ( .D(\row1_buffer[172][3] ), .CK(clk), .Q(
        \row1_buffer[171][3] ) );
  DFFQXL \row1_buffer_reg[170][3]  ( .D(\row1_buffer[171][3] ), .CK(clk), .Q(
        \row1_buffer[170][3] ) );
  DFFQXL \row1_buffer_reg[169][3]  ( .D(\row1_buffer[170][3] ), .CK(clk), .Q(
        \row1_buffer[169][3] ) );
  DFFQXL \row1_buffer_reg[168][3]  ( .D(\row1_buffer[169][3] ), .CK(clk), .Q(
        \row1_buffer[168][3] ) );
  DFFQXL \row1_buffer_reg[167][3]  ( .D(\row1_buffer[168][3] ), .CK(clk), .Q(
        \row1_buffer[167][3] ) );
  DFFQXL \row1_buffer_reg[166][3]  ( .D(\row1_buffer[167][3] ), .CK(clk), .Q(
        \row1_buffer[166][3] ) );
  DFFQXL \row1_buffer_reg[165][3]  ( .D(\row1_buffer[166][3] ), .CK(clk), .Q(
        \row1_buffer[165][3] ) );
  DFFQXL \row1_buffer_reg[164][3]  ( .D(\row1_buffer[165][3] ), .CK(clk), .Q(
        \row1_buffer[164][3] ) );
  DFFQXL \row1_buffer_reg[163][3]  ( .D(\row1_buffer[164][3] ), .CK(clk), .Q(
        \row1_buffer[163][3] ) );
  DFFQXL \row1_buffer_reg[162][3]  ( .D(\row1_buffer[163][3] ), .CK(clk), .Q(
        \row1_buffer[162][3] ) );
  DFFQXL \row1_buffer_reg[161][3]  ( .D(\row1_buffer[162][3] ), .CK(clk), .Q(
        \row1_buffer[161][3] ) );
  DFFQXL \row1_buffer_reg[160][3]  ( .D(\row1_buffer[161][3] ), .CK(clk), .Q(
        \row1_buffer[160][3] ) );
  DFFQXL \row1_buffer_reg[159][3]  ( .D(\row1_buffer[160][3] ), .CK(clk), .Q(
        \row1_buffer[159][3] ) );
  DFFQXL \row1_buffer_reg[158][3]  ( .D(\row1_buffer[159][3] ), .CK(clk), .Q(
        \row1_buffer[158][3] ) );
  DFFQXL \row1_buffer_reg[157][3]  ( .D(\row1_buffer[158][3] ), .CK(clk), .Q(
        \row1_buffer[157][3] ) );
  DFFQXL \row1_buffer_reg[156][3]  ( .D(\row1_buffer[157][3] ), .CK(clk), .Q(
        \row1_buffer[156][3] ) );
  DFFQXL \row1_buffer_reg[155][3]  ( .D(\row1_buffer[156][3] ), .CK(clk), .Q(
        \row1_buffer[155][3] ) );
  DFFQXL \row1_buffer_reg[154][3]  ( .D(\row1_buffer[155][3] ), .CK(clk), .Q(
        \row1_buffer[154][3] ) );
  DFFQXL \row1_buffer_reg[153][3]  ( .D(\row1_buffer[154][3] ), .CK(clk), .Q(
        \row1_buffer[153][3] ) );
  DFFQXL \row1_buffer_reg[152][3]  ( .D(\row1_buffer[153][3] ), .CK(clk), .Q(
        \row1_buffer[152][3] ) );
  DFFQXL \row1_buffer_reg[151][3]  ( .D(\row1_buffer[152][3] ), .CK(clk), .Q(
        \row1_buffer[151][3] ) );
  DFFQXL \row1_buffer_reg[150][3]  ( .D(\row1_buffer[151][3] ), .CK(clk), .Q(
        \row1_buffer[150][3] ) );
  DFFQXL \row1_buffer_reg[149][3]  ( .D(\row1_buffer[150][3] ), .CK(clk), .Q(
        \row1_buffer[149][3] ) );
  DFFQXL \row1_buffer_reg[148][3]  ( .D(\row1_buffer[149][3] ), .CK(clk), .Q(
        \row1_buffer[148][3] ) );
  DFFQXL \row1_buffer_reg[147][3]  ( .D(\row1_buffer[148][3] ), .CK(clk), .Q(
        \row1_buffer[147][3] ) );
  DFFQXL \row1_buffer_reg[146][3]  ( .D(\row1_buffer[147][3] ), .CK(clk), .Q(
        \row1_buffer[146][3] ) );
  DFFQXL \row1_buffer_reg[145][3]  ( .D(\row1_buffer[146][3] ), .CK(clk), .Q(
        \row1_buffer[145][3] ) );
  DFFQXL \row1_buffer_reg[144][3]  ( .D(\row1_buffer[145][3] ), .CK(clk), .Q(
        \row1_buffer[144][3] ) );
  DFFQXL \row1_buffer_reg[143][3]  ( .D(\row1_buffer[144][3] ), .CK(clk), .Q(
        \row1_buffer[143][3] ) );
  DFFQXL \row1_buffer_reg[142][3]  ( .D(\row1_buffer[143][3] ), .CK(clk), .Q(
        \row1_buffer[142][3] ) );
  DFFQXL \row1_buffer_reg[141][3]  ( .D(\row1_buffer[142][3] ), .CK(clk), .Q(
        \row1_buffer[141][3] ) );
  DFFQXL \row1_buffer_reg[140][3]  ( .D(\row1_buffer[141][3] ), .CK(clk), .Q(
        \row1_buffer[140][3] ) );
  DFFQXL \row1_buffer_reg[139][3]  ( .D(\row1_buffer[140][3] ), .CK(clk), .Q(
        \row1_buffer[139][3] ) );
  DFFQXL \row1_buffer_reg[138][3]  ( .D(\row1_buffer[139][3] ), .CK(clk), .Q(
        \row1_buffer[138][3] ) );
  DFFQXL \row1_buffer_reg[137][3]  ( .D(\row1_buffer[138][3] ), .CK(clk), .Q(
        \row1_buffer[137][3] ) );
  DFFQXL \row1_buffer_reg[136][3]  ( .D(\row1_buffer[137][3] ), .CK(clk), .Q(
        \row1_buffer[136][3] ) );
  DFFQXL \row1_buffer_reg[135][3]  ( .D(\row1_buffer[136][3] ), .CK(clk), .Q(
        \row1_buffer[135][3] ) );
  DFFQXL \row1_buffer_reg[134][3]  ( .D(\row1_buffer[135][3] ), .CK(clk), .Q(
        \row1_buffer[134][3] ) );
  DFFQXL \row1_buffer_reg[133][3]  ( .D(\row1_buffer[134][3] ), .CK(clk), .Q(
        \row1_buffer[133][3] ) );
  DFFQXL \row1_buffer_reg[132][3]  ( .D(\row1_buffer[133][3] ), .CK(clk), .Q(
        \row1_buffer[132][3] ) );
  DFFQXL \row1_buffer_reg[131][3]  ( .D(\row1_buffer[132][3] ), .CK(clk), .Q(
        \row1_buffer[131][3] ) );
  DFFQXL \row1_buffer_reg[130][3]  ( .D(\row1_buffer[131][3] ), .CK(clk), .Q(
        \row1_buffer[130][3] ) );
  DFFQXL \row1_buffer_reg[129][3]  ( .D(\row1_buffer[130][3] ), .CK(clk), .Q(
        \row1_buffer[129][3] ) );
  DFFQXL \row1_buffer_reg[128][3]  ( .D(\row1_buffer[129][3] ), .CK(clk), .Q(
        \row1_buffer[128][3] ) );
  DFFQXL \row1_buffer_reg[127][3]  ( .D(\row1_buffer[128][3] ), .CK(clk), .Q(
        \row1_buffer[127][3] ) );
  DFFQXL \row1_buffer_reg[126][3]  ( .D(\row1_buffer[127][3] ), .CK(clk), .Q(
        \row1_buffer[126][3] ) );
  DFFQXL \row1_buffer_reg[125][3]  ( .D(\row1_buffer[126][3] ), .CK(clk), .Q(
        \row1_buffer[125][3] ) );
  DFFQXL \row1_buffer_reg[124][3]  ( .D(\row1_buffer[125][3] ), .CK(clk), .Q(
        \row1_buffer[124][3] ) );
  DFFQXL \row1_buffer_reg[123][3]  ( .D(\row1_buffer[124][3] ), .CK(clk), .Q(
        \row1_buffer[123][3] ) );
  DFFQXL \row1_buffer_reg[122][3]  ( .D(\row1_buffer[123][3] ), .CK(clk), .Q(
        \row1_buffer[122][3] ) );
  DFFQXL \row1_buffer_reg[121][3]  ( .D(\row1_buffer[122][3] ), .CK(clk), .Q(
        \row1_buffer[121][3] ) );
  DFFQXL \row1_buffer_reg[120][3]  ( .D(\row1_buffer[121][3] ), .CK(clk), .Q(
        \row1_buffer[120][3] ) );
  DFFQXL \row1_buffer_reg[119][3]  ( .D(\row1_buffer[120][3] ), .CK(clk), .Q(
        \row1_buffer[119][3] ) );
  DFFQXL \row1_buffer_reg[118][3]  ( .D(\row1_buffer[119][3] ), .CK(clk), .Q(
        \row1_buffer[118][3] ) );
  DFFQXL \row1_buffer_reg[117][3]  ( .D(\row1_buffer[118][3] ), .CK(clk), .Q(
        \row1_buffer[117][3] ) );
  DFFQXL \row1_buffer_reg[116][3]  ( .D(\row1_buffer[117][3] ), .CK(clk), .Q(
        \row1_buffer[116][3] ) );
  DFFQXL \row1_buffer_reg[115][3]  ( .D(\row1_buffer[116][3] ), .CK(clk), .Q(
        \row1_buffer[115][3] ) );
  DFFQXL \row1_buffer_reg[114][3]  ( .D(\row1_buffer[115][3] ), .CK(clk), .Q(
        \row1_buffer[114][3] ) );
  DFFQXL \row1_buffer_reg[113][3]  ( .D(\row1_buffer[114][3] ), .CK(clk), .Q(
        \row1_buffer[113][3] ) );
  DFFQXL \row1_buffer_reg[112][3]  ( .D(\row1_buffer[113][3] ), .CK(clk), .Q(
        \row1_buffer[112][3] ) );
  DFFQXL \row1_buffer_reg[111][3]  ( .D(\row1_buffer[112][3] ), .CK(clk), .Q(
        \row1_buffer[111][3] ) );
  DFFQXL \row1_buffer_reg[110][3]  ( .D(\row1_buffer[111][3] ), .CK(clk), .Q(
        \row1_buffer[110][3] ) );
  DFFQXL \row1_buffer_reg[109][3]  ( .D(\row1_buffer[110][3] ), .CK(clk), .Q(
        \row1_buffer[109][3] ) );
  DFFQXL \row1_buffer_reg[108][3]  ( .D(\row1_buffer[109][3] ), .CK(clk), .Q(
        \row1_buffer[108][3] ) );
  DFFQXL \row1_buffer_reg[107][3]  ( .D(\row1_buffer[108][3] ), .CK(clk), .Q(
        \row1_buffer[107][3] ) );
  DFFQXL \row1_buffer_reg[106][3]  ( .D(\row1_buffer[107][3] ), .CK(clk), .Q(
        \row1_buffer[106][3] ) );
  DFFQXL \row1_buffer_reg[105][3]  ( .D(\row1_buffer[106][3] ), .CK(clk), .Q(
        \row1_buffer[105][3] ) );
  DFFQXL \row1_buffer_reg[104][3]  ( .D(\row1_buffer[105][3] ), .CK(clk), .Q(
        \row1_buffer[104][3] ) );
  DFFQXL \row1_buffer_reg[103][3]  ( .D(\row1_buffer[104][3] ), .CK(clk), .Q(
        \row1_buffer[103][3] ) );
  DFFQXL \row1_buffer_reg[102][3]  ( .D(\row1_buffer[103][3] ), .CK(clk), .Q(
        \row1_buffer[102][3] ) );
  DFFQXL \row1_buffer_reg[101][3]  ( .D(\row1_buffer[102][3] ), .CK(clk), .Q(
        \row1_buffer[101][3] ) );
  DFFQXL \row1_buffer_reg[100][3]  ( .D(\row1_buffer[101][3] ), .CK(clk), .Q(
        \row1_buffer[100][3] ) );
  DFFQXL \row1_buffer_reg[99][3]  ( .D(\row1_buffer[100][3] ), .CK(clk), .Q(
        \row1_buffer[99][3] ) );
  DFFQXL \row1_buffer_reg[98][3]  ( .D(\row1_buffer[99][3] ), .CK(clk), .Q(
        \row1_buffer[98][3] ) );
  DFFQXL \row1_buffer_reg[97][3]  ( .D(\row1_buffer[98][3] ), .CK(clk), .Q(
        \row1_buffer[97][3] ) );
  DFFQXL \row1_buffer_reg[96][3]  ( .D(\row1_buffer[97][3] ), .CK(clk), .Q(
        \row1_buffer[96][3] ) );
  DFFQXL \row1_buffer_reg[95][3]  ( .D(\row1_buffer[96][3] ), .CK(clk), .Q(
        \row1_buffer[95][3] ) );
  DFFQXL \row1_buffer_reg[94][3]  ( .D(\row1_buffer[95][3] ), .CK(clk), .Q(
        \row1_buffer[94][3] ) );
  DFFQXL \row1_buffer_reg[93][3]  ( .D(\row1_buffer[94][3] ), .CK(clk), .Q(
        \row1_buffer[93][3] ) );
  DFFQXL \row1_buffer_reg[92][3]  ( .D(\row1_buffer[93][3] ), .CK(clk), .Q(
        \row1_buffer[92][3] ) );
  DFFQXL \row1_buffer_reg[91][3]  ( .D(\row1_buffer[92][3] ), .CK(clk), .Q(
        \row1_buffer[91][3] ) );
  DFFQXL \row1_buffer_reg[90][3]  ( .D(\row1_buffer[91][3] ), .CK(clk), .Q(
        \row1_buffer[90][3] ) );
  DFFQXL \row1_buffer_reg[89][3]  ( .D(\row1_buffer[90][3] ), .CK(clk), .Q(
        \row1_buffer[89][3] ) );
  DFFQXL \row1_buffer_reg[88][3]  ( .D(\row1_buffer[89][3] ), .CK(clk), .Q(
        \row1_buffer[88][3] ) );
  DFFQXL \row1_buffer_reg[87][3]  ( .D(\row1_buffer[88][3] ), .CK(clk), .Q(
        \row1_buffer[87][3] ) );
  DFFQXL \row1_buffer_reg[86][3]  ( .D(\row1_buffer[87][3] ), .CK(clk), .Q(
        \row1_buffer[86][3] ) );
  DFFQXL \row1_buffer_reg[85][3]  ( .D(\row1_buffer[86][3] ), .CK(clk), .Q(
        \row1_buffer[85][3] ) );
  DFFQXL \row1_buffer_reg[84][3]  ( .D(\row1_buffer[85][3] ), .CK(clk), .Q(
        \row1_buffer[84][3] ) );
  DFFQXL \row1_buffer_reg[83][3]  ( .D(\row1_buffer[84][3] ), .CK(clk), .Q(
        \row1_buffer[83][3] ) );
  DFFQXL \row1_buffer_reg[82][3]  ( .D(\row1_buffer[83][3] ), .CK(clk), .Q(
        \row1_buffer[82][3] ) );
  DFFQXL \row1_buffer_reg[81][3]  ( .D(\row1_buffer[82][3] ), .CK(clk), .Q(
        \row1_buffer[81][3] ) );
  DFFQXL \row1_buffer_reg[80][3]  ( .D(\row1_buffer[81][3] ), .CK(clk), .Q(
        \row1_buffer[80][3] ) );
  DFFQXL \row1_buffer_reg[79][3]  ( .D(\row1_buffer[80][3] ), .CK(clk), .Q(
        \row1_buffer[79][3] ) );
  DFFQXL \row1_buffer_reg[78][3]  ( .D(\row1_buffer[79][3] ), .CK(clk), .Q(
        \row1_buffer[78][3] ) );
  DFFQXL \row1_buffer_reg[77][3]  ( .D(\row1_buffer[78][3] ), .CK(clk), .Q(
        \row1_buffer[77][3] ) );
  DFFQXL \row1_buffer_reg[76][3]  ( .D(\row1_buffer[77][3] ), .CK(clk), .Q(
        \row1_buffer[76][3] ) );
  DFFQXL \row1_buffer_reg[75][3]  ( .D(\row1_buffer[76][3] ), .CK(clk), .Q(
        \row1_buffer[75][3] ) );
  DFFQXL \row1_buffer_reg[74][3]  ( .D(\row1_buffer[75][3] ), .CK(clk), .Q(
        \row1_buffer[74][3] ) );
  DFFQXL \row1_buffer_reg[73][3]  ( .D(\row1_buffer[74][3] ), .CK(clk), .Q(
        \row1_buffer[73][3] ) );
  DFFQXL \row1_buffer_reg[72][3]  ( .D(\row1_buffer[73][3] ), .CK(clk), .Q(
        \row1_buffer[72][3] ) );
  DFFQXL \row1_buffer_reg[71][3]  ( .D(\row1_buffer[72][3] ), .CK(clk), .Q(
        \row1_buffer[71][3] ) );
  DFFQXL \row1_buffer_reg[70][3]  ( .D(\row1_buffer[71][3] ), .CK(clk), .Q(
        \row1_buffer[70][3] ) );
  DFFQXL \row1_buffer_reg[69][3]  ( .D(\row1_buffer[70][3] ), .CK(clk), .Q(
        \row1_buffer[69][3] ) );
  DFFQXL \row1_buffer_reg[68][3]  ( .D(\row1_buffer[69][3] ), .CK(clk), .Q(
        \row1_buffer[68][3] ) );
  DFFQXL \row1_buffer_reg[67][3]  ( .D(\row1_buffer[68][3] ), .CK(clk), .Q(
        \row1_buffer[67][3] ) );
  DFFQXL \row1_buffer_reg[66][3]  ( .D(\row1_buffer[67][3] ), .CK(clk), .Q(
        \row1_buffer[66][3] ) );
  DFFQXL \row1_buffer_reg[65][3]  ( .D(\row1_buffer[66][3] ), .CK(clk), .Q(
        \row1_buffer[65][3] ) );
  DFFQXL \row1_buffer_reg[64][3]  ( .D(\row1_buffer[65][3] ), .CK(clk), .Q(
        \row1_buffer[64][3] ) );
  DFFQXL \row1_buffer_reg[63][3]  ( .D(\row1_buffer[64][3] ), .CK(clk), .Q(
        \row1_buffer[63][3] ) );
  DFFQXL \row1_buffer_reg[62][3]  ( .D(\row1_buffer[63][3] ), .CK(clk), .Q(
        \row1_buffer[62][3] ) );
  DFFQXL \row1_buffer_reg[61][3]  ( .D(\row1_buffer[62][3] ), .CK(clk), .Q(
        \row1_buffer[61][3] ) );
  DFFQXL \row1_buffer_reg[60][3]  ( .D(\row1_buffer[61][3] ), .CK(clk), .Q(
        \row1_buffer[60][3] ) );
  DFFQXL \row1_buffer_reg[59][3]  ( .D(\row1_buffer[60][3] ), .CK(clk), .Q(
        \row1_buffer[59][3] ) );
  DFFQXL \row1_buffer_reg[58][3]  ( .D(\row1_buffer[59][3] ), .CK(clk), .Q(
        \row1_buffer[58][3] ) );
  DFFQXL \row1_buffer_reg[57][3]  ( .D(\row1_buffer[58][3] ), .CK(clk), .Q(
        \row1_buffer[57][3] ) );
  DFFQXL \row1_buffer_reg[56][3]  ( .D(\row1_buffer[57][3] ), .CK(clk), .Q(
        \row1_buffer[56][3] ) );
  DFFQXL \row1_buffer_reg[55][3]  ( .D(\row1_buffer[56][3] ), .CK(clk), .Q(
        \row1_buffer[55][3] ) );
  DFFQXL \row1_buffer_reg[54][3]  ( .D(\row1_buffer[55][3] ), .CK(clk), .Q(
        \row1_buffer[54][3] ) );
  DFFQXL \row1_buffer_reg[53][3]  ( .D(\row1_buffer[54][3] ), .CK(clk), .Q(
        \row1_buffer[53][3] ) );
  DFFQXL \row1_buffer_reg[52][3]  ( .D(\row1_buffer[53][3] ), .CK(clk), .Q(
        \row1_buffer[52][3] ) );
  DFFQXL \row1_buffer_reg[51][3]  ( .D(\row1_buffer[52][3] ), .CK(clk), .Q(
        \row1_buffer[51][3] ) );
  DFFQXL \row1_buffer_reg[50][3]  ( .D(\row1_buffer[51][3] ), .CK(clk), .Q(
        \row1_buffer[50][3] ) );
  DFFQXL \row1_buffer_reg[49][3]  ( .D(\row1_buffer[50][3] ), .CK(clk), .Q(
        \row1_buffer[49][3] ) );
  DFFQXL \row1_buffer_reg[48][3]  ( .D(\row1_buffer[49][3] ), .CK(clk), .Q(
        \row1_buffer[48][3] ) );
  DFFQXL \row1_buffer_reg[47][3]  ( .D(\row1_buffer[48][3] ), .CK(clk), .Q(
        \row1_buffer[47][3] ) );
  DFFQXL \row1_buffer_reg[46][3]  ( .D(\row1_buffer[47][3] ), .CK(clk), .Q(
        \row1_buffer[46][3] ) );
  DFFQXL \row1_buffer_reg[45][3]  ( .D(\row1_buffer[46][3] ), .CK(clk), .Q(
        \row1_buffer[45][3] ) );
  DFFQXL \row1_buffer_reg[44][3]  ( .D(\row1_buffer[45][3] ), .CK(clk), .Q(
        \row1_buffer[44][3] ) );
  DFFQXL \row1_buffer_reg[43][3]  ( .D(\row1_buffer[44][3] ), .CK(clk), .Q(
        \row1_buffer[43][3] ) );
  DFFQXL \row1_buffer_reg[42][3]  ( .D(\row1_buffer[43][3] ), .CK(clk), .Q(
        \row1_buffer[42][3] ) );
  DFFQXL \row1_buffer_reg[41][3]  ( .D(\row1_buffer[42][3] ), .CK(clk), .Q(
        \row1_buffer[41][3] ) );
  DFFQXL \row1_buffer_reg[40][3]  ( .D(\row1_buffer[41][3] ), .CK(clk), .Q(
        \row1_buffer[40][3] ) );
  DFFQXL \row1_buffer_reg[39][3]  ( .D(\row1_buffer[40][3] ), .CK(clk), .Q(
        \row1_buffer[39][3] ) );
  DFFQXL \row1_buffer_reg[38][3]  ( .D(\row1_buffer[39][3] ), .CK(clk), .Q(
        \row1_buffer[38][3] ) );
  DFFQXL \row1_buffer_reg[37][3]  ( .D(\row1_buffer[38][3] ), .CK(clk), .Q(
        \row1_buffer[37][3] ) );
  DFFQXL \row1_buffer_reg[36][3]  ( .D(\row1_buffer[37][3] ), .CK(clk), .Q(
        \row1_buffer[36][3] ) );
  DFFQXL \row1_buffer_reg[35][3]  ( .D(\row1_buffer[36][3] ), .CK(clk), .Q(
        \row1_buffer[35][3] ) );
  DFFQXL \row1_buffer_reg[34][3]  ( .D(\row1_buffer[35][3] ), .CK(clk), .Q(
        \row1_buffer[34][3] ) );
  DFFQXL \row1_buffer_reg[33][3]  ( .D(\row1_buffer[34][3] ), .CK(clk), .Q(
        \row1_buffer[33][3] ) );
  DFFQXL \row1_buffer_reg[32][3]  ( .D(\row1_buffer[33][3] ), .CK(clk), .Q(
        \row1_buffer[32][3] ) );
  DFFQXL \row1_buffer_reg[31][3]  ( .D(\row1_buffer[32][3] ), .CK(clk), .Q(
        \row1_buffer[31][3] ) );
  DFFQXL \row1_buffer_reg[30][3]  ( .D(\row1_buffer[31][3] ), .CK(clk), .Q(
        \row1_buffer[30][3] ) );
  DFFQXL \row1_buffer_reg[29][3]  ( .D(\row1_buffer[30][3] ), .CK(clk), .Q(
        \row1_buffer[29][3] ) );
  DFFQXL \row1_buffer_reg[28][3]  ( .D(\row1_buffer[29][3] ), .CK(clk), .Q(
        \row1_buffer[28][3] ) );
  DFFQXL \row1_buffer_reg[27][3]  ( .D(\row1_buffer[28][3] ), .CK(clk), .Q(
        \row1_buffer[27][3] ) );
  DFFQXL \row1_buffer_reg[26][3]  ( .D(\row1_buffer[27][3] ), .CK(clk), .Q(
        \row1_buffer[26][3] ) );
  DFFQXL \row1_buffer_reg[25][3]  ( .D(\row1_buffer[26][3] ), .CK(clk), .Q(
        \row1_buffer[25][3] ) );
  DFFQXL \row1_buffer_reg[24][3]  ( .D(\row1_buffer[25][3] ), .CK(clk), .Q(
        \row1_buffer[24][3] ) );
  DFFQXL \row1_buffer_reg[23][3]  ( .D(\row1_buffer[24][3] ), .CK(clk), .Q(
        \row1_buffer[23][3] ) );
  DFFQXL \row1_buffer_reg[22][3]  ( .D(\row1_buffer[23][3] ), .CK(clk), .Q(
        \row1_buffer[22][3] ) );
  DFFQXL \row1_buffer_reg[21][3]  ( .D(\row1_buffer[22][3] ), .CK(clk), .Q(
        \row1_buffer[21][3] ) );
  DFFQXL \row1_buffer_reg[20][3]  ( .D(\row1_buffer[21][3] ), .CK(clk), .Q(
        \row1_buffer[20][3] ) );
  DFFQXL \row1_buffer_reg[19][3]  ( .D(\row1_buffer[20][3] ), .CK(clk), .Q(
        \row1_buffer[19][3] ) );
  DFFQXL \row1_buffer_reg[18][3]  ( .D(\row1_buffer[19][3] ), .CK(clk), .Q(
        \row1_buffer[18][3] ) );
  DFFQXL \row1_buffer_reg[17][3]  ( .D(\row1_buffer[18][3] ), .CK(clk), .Q(
        \row1_buffer[17][3] ) );
  DFFQXL \row1_buffer_reg[16][3]  ( .D(\row1_buffer[17][3] ), .CK(clk), .Q(
        \row1_buffer[16][3] ) );
  DFFQXL \row1_buffer_reg[15][3]  ( .D(\row1_buffer[16][3] ), .CK(clk), .Q(
        \row1_buffer[15][3] ) );
  DFFQXL \row1_buffer_reg[14][3]  ( .D(\row1_buffer[15][3] ), .CK(clk), .Q(
        \row1_buffer[14][3] ) );
  DFFQXL \row1_buffer_reg[13][3]  ( .D(\row1_buffer[14][3] ), .CK(clk), .Q(
        \row1_buffer[13][3] ) );
  DFFQXL \row1_buffer_reg[12][3]  ( .D(\row1_buffer[13][3] ), .CK(clk), .Q(
        \row1_buffer[12][3] ) );
  DFFQXL \row1_buffer_reg[11][3]  ( .D(\row1_buffer[12][3] ), .CK(clk), .Q(
        \row1_buffer[11][3] ) );
  DFFQXL \row1_buffer_reg[10][3]  ( .D(\row1_buffer[11][3] ), .CK(clk), .Q(
        \row1_buffer[10][3] ) );
  DFFQXL \row1_buffer_reg[9][3]  ( .D(\row1_buffer[10][3] ), .CK(clk), .Q(
        \row1_buffer[9][3] ) );
  DFFQXL \row1_buffer_reg[8][3]  ( .D(\row1_buffer[9][3] ), .CK(clk), .Q(
        \row1_buffer[8][3] ) );
  DFFQXL \row1_buffer_reg[7][3]  ( .D(\row1_buffer[8][3] ), .CK(clk), .Q(
        \row1_buffer[7][3] ) );
  DFFQXL \row1_buffer_reg[6][3]  ( .D(\row1_buffer[7][3] ), .CK(clk), .Q(
        \row1_buffer[6][3] ) );
  DFFQXL \row1_buffer_reg[5][3]  ( .D(\row1_buffer[6][3] ), .CK(clk), .Q(
        \row1_buffer[5][3] ) );
  DFFQXL \row1_buffer_reg[4][3]  ( .D(\row1_buffer[5][3] ), .CK(clk), .Q(
        \row1_buffer[4][3] ) );
  DFFQXL \row1_buffer_reg[3][3]  ( .D(\row1_buffer[4][3] ), .CK(clk), .Q(
        \row1_buffer[3][3] ) );
  DFFQXL \row1_buffer_reg[0][3]  ( .D(\row1_buffer[1][3] ), .CK(clk), .Q(
        \row1_buffer[0][3] ) );
  DFFQXL \row2_buffer_reg[225][2]  ( .D(\row3_buffer[0][2] ), .CK(clk), .Q(
        \row2_buffer[225][2] ) );
  DFFQXL \row2_buffer_reg[224][2]  ( .D(\row2_buffer[225][2] ), .CK(clk), .Q(
        \row2_buffer[224][2] ) );
  DFFQXL \row2_buffer_reg[223][2]  ( .D(\row2_buffer[224][2] ), .CK(clk), .Q(
        \row2_buffer[223][2] ) );
  DFFQXL \row2_buffer_reg[222][2]  ( .D(\row2_buffer[223][2] ), .CK(clk), .Q(
        \row2_buffer[222][2] ) );
  DFFQXL \row2_buffer_reg[221][2]  ( .D(\row2_buffer[222][2] ), .CK(clk), .Q(
        \row2_buffer[221][2] ) );
  DFFQXL \row2_buffer_reg[220][2]  ( .D(\row2_buffer[221][2] ), .CK(clk), .Q(
        \row2_buffer[220][2] ) );
  DFFQXL \row2_buffer_reg[219][2]  ( .D(\row2_buffer[220][2] ), .CK(clk), .Q(
        \row2_buffer[219][2] ) );
  DFFQXL \row2_buffer_reg[218][2]  ( .D(\row2_buffer[219][2] ), .CK(clk), .Q(
        \row2_buffer[218][2] ) );
  DFFQXL \row2_buffer_reg[217][2]  ( .D(\row2_buffer[218][2] ), .CK(clk), .Q(
        \row2_buffer[217][2] ) );
  DFFQXL \row2_buffer_reg[216][2]  ( .D(\row2_buffer[217][2] ), .CK(clk), .Q(
        \row2_buffer[216][2] ) );
  DFFQXL \row2_buffer_reg[215][2]  ( .D(\row2_buffer[216][2] ), .CK(clk), .Q(
        \row2_buffer[215][2] ) );
  DFFQXL \row2_buffer_reg[214][2]  ( .D(\row2_buffer[215][2] ), .CK(clk), .Q(
        \row2_buffer[214][2] ) );
  DFFQXL \row2_buffer_reg[213][2]  ( .D(\row2_buffer[214][2] ), .CK(clk), .Q(
        \row2_buffer[213][2] ) );
  DFFQXL \row2_buffer_reg[212][2]  ( .D(\row2_buffer[213][2] ), .CK(clk), .Q(
        \row2_buffer[212][2] ) );
  DFFQXL \row2_buffer_reg[211][2]  ( .D(\row2_buffer[212][2] ), .CK(clk), .Q(
        \row2_buffer[211][2] ) );
  DFFQXL \row2_buffer_reg[210][2]  ( .D(\row2_buffer[211][2] ), .CK(clk), .Q(
        \row2_buffer[210][2] ) );
  DFFQXL \row2_buffer_reg[209][2]  ( .D(\row2_buffer[210][2] ), .CK(clk), .Q(
        \row2_buffer[209][2] ) );
  DFFQXL \row2_buffer_reg[208][2]  ( .D(\row2_buffer[209][2] ), .CK(clk), .Q(
        \row2_buffer[208][2] ) );
  DFFQXL \row2_buffer_reg[207][2]  ( .D(\row2_buffer[208][2] ), .CK(clk), .Q(
        \row2_buffer[207][2] ) );
  DFFQXL \row2_buffer_reg[206][2]  ( .D(\row2_buffer[207][2] ), .CK(clk), .Q(
        \row2_buffer[206][2] ) );
  DFFQXL \row2_buffer_reg[205][2]  ( .D(\row2_buffer[206][2] ), .CK(clk), .Q(
        \row2_buffer[205][2] ) );
  DFFQXL \row2_buffer_reg[204][2]  ( .D(\row2_buffer[205][2] ), .CK(clk), .Q(
        \row2_buffer[204][2] ) );
  DFFQXL \row2_buffer_reg[203][2]  ( .D(\row2_buffer[204][2] ), .CK(clk), .Q(
        \row2_buffer[203][2] ) );
  DFFQXL \row2_buffer_reg[202][2]  ( .D(\row2_buffer[203][2] ), .CK(clk), .Q(
        \row2_buffer[202][2] ) );
  DFFQXL \row2_buffer_reg[201][2]  ( .D(\row2_buffer[202][2] ), .CK(clk), .Q(
        \row2_buffer[201][2] ) );
  DFFQXL \row2_buffer_reg[200][2]  ( .D(\row2_buffer[201][2] ), .CK(clk), .Q(
        \row2_buffer[200][2] ) );
  DFFQXL \row2_buffer_reg[199][2]  ( .D(\row2_buffer[200][2] ), .CK(clk), .Q(
        \row2_buffer[199][2] ) );
  DFFQXL \row2_buffer_reg[198][2]  ( .D(\row2_buffer[199][2] ), .CK(clk), .Q(
        \row2_buffer[198][2] ) );
  DFFQXL \row2_buffer_reg[197][2]  ( .D(\row2_buffer[198][2] ), .CK(clk), .Q(
        \row2_buffer[197][2] ) );
  DFFQXL \row2_buffer_reg[196][2]  ( .D(\row2_buffer[197][2] ), .CK(clk), .Q(
        \row2_buffer[196][2] ) );
  DFFQXL \row2_buffer_reg[195][2]  ( .D(\row2_buffer[196][2] ), .CK(clk), .Q(
        \row2_buffer[195][2] ) );
  DFFQXL \row2_buffer_reg[194][2]  ( .D(\row2_buffer[195][2] ), .CK(clk), .Q(
        \row2_buffer[194][2] ) );
  DFFQXL \row2_buffer_reg[193][2]  ( .D(\row2_buffer[194][2] ), .CK(clk), .Q(
        \row2_buffer[193][2] ) );
  DFFQXL \row2_buffer_reg[192][2]  ( .D(\row2_buffer[193][2] ), .CK(clk), .Q(
        \row2_buffer[192][2] ) );
  DFFQXL \row2_buffer_reg[191][2]  ( .D(\row2_buffer[192][2] ), .CK(clk), .Q(
        \row2_buffer[191][2] ) );
  DFFQXL \row2_buffer_reg[190][2]  ( .D(\row2_buffer[191][2] ), .CK(clk), .Q(
        \row2_buffer[190][2] ) );
  DFFQXL \row2_buffer_reg[189][2]  ( .D(\row2_buffer[190][2] ), .CK(clk), .Q(
        \row2_buffer[189][2] ) );
  DFFQXL \row2_buffer_reg[188][2]  ( .D(\row2_buffer[189][2] ), .CK(clk), .Q(
        \row2_buffer[188][2] ) );
  DFFQXL \row2_buffer_reg[187][2]  ( .D(\row2_buffer[188][2] ), .CK(clk), .Q(
        \row2_buffer[187][2] ) );
  DFFQXL \row2_buffer_reg[186][2]  ( .D(\row2_buffer[187][2] ), .CK(clk), .Q(
        \row2_buffer[186][2] ) );
  DFFQXL \row2_buffer_reg[185][2]  ( .D(\row2_buffer[186][2] ), .CK(clk), .Q(
        \row2_buffer[185][2] ) );
  DFFQXL \row2_buffer_reg[184][2]  ( .D(\row2_buffer[185][2] ), .CK(clk), .Q(
        \row2_buffer[184][2] ) );
  DFFQXL \row2_buffer_reg[183][2]  ( .D(\row2_buffer[184][2] ), .CK(clk), .Q(
        \row2_buffer[183][2] ) );
  DFFQXL \row2_buffer_reg[182][2]  ( .D(\row2_buffer[183][2] ), .CK(clk), .Q(
        \row2_buffer[182][2] ) );
  DFFQXL \row2_buffer_reg[181][2]  ( .D(\row2_buffer[182][2] ), .CK(clk), .Q(
        \row2_buffer[181][2] ) );
  DFFQXL \row2_buffer_reg[180][2]  ( .D(\row2_buffer[181][2] ), .CK(clk), .Q(
        \row2_buffer[180][2] ) );
  DFFQXL \row2_buffer_reg[179][2]  ( .D(\row2_buffer[180][2] ), .CK(clk), .Q(
        \row2_buffer[179][2] ) );
  DFFQXL \row2_buffer_reg[178][2]  ( .D(\row2_buffer[179][2] ), .CK(clk), .Q(
        \row2_buffer[178][2] ) );
  DFFQXL \row2_buffer_reg[177][2]  ( .D(\row2_buffer[178][2] ), .CK(clk), .Q(
        \row2_buffer[177][2] ) );
  DFFQXL \row2_buffer_reg[176][2]  ( .D(\row2_buffer[177][2] ), .CK(clk), .Q(
        \row2_buffer[176][2] ) );
  DFFQXL \row2_buffer_reg[175][2]  ( .D(\row2_buffer[176][2] ), .CK(clk), .Q(
        \row2_buffer[175][2] ) );
  DFFQXL \row2_buffer_reg[174][2]  ( .D(\row2_buffer[175][2] ), .CK(clk), .Q(
        \row2_buffer[174][2] ) );
  DFFQXL \row2_buffer_reg[173][2]  ( .D(\row2_buffer[174][2] ), .CK(clk), .Q(
        \row2_buffer[173][2] ) );
  DFFQXL \row2_buffer_reg[172][2]  ( .D(\row2_buffer[173][2] ), .CK(clk), .Q(
        \row2_buffer[172][2] ) );
  DFFQXL \row2_buffer_reg[171][2]  ( .D(\row2_buffer[172][2] ), .CK(clk), .Q(
        \row2_buffer[171][2] ) );
  DFFQXL \row2_buffer_reg[170][2]  ( .D(\row2_buffer[171][2] ), .CK(clk), .Q(
        \row2_buffer[170][2] ) );
  DFFQXL \row2_buffer_reg[169][2]  ( .D(\row2_buffer[170][2] ), .CK(clk), .Q(
        \row2_buffer[169][2] ) );
  DFFQXL \row2_buffer_reg[168][2]  ( .D(\row2_buffer[169][2] ), .CK(clk), .Q(
        \row2_buffer[168][2] ) );
  DFFQXL \row2_buffer_reg[167][2]  ( .D(\row2_buffer[168][2] ), .CK(clk), .Q(
        \row2_buffer[167][2] ) );
  DFFQXL \row2_buffer_reg[166][2]  ( .D(\row2_buffer[167][2] ), .CK(clk), .Q(
        \row2_buffer[166][2] ) );
  DFFQXL \row2_buffer_reg[165][2]  ( .D(\row2_buffer[166][2] ), .CK(clk), .Q(
        \row2_buffer[165][2] ) );
  DFFQXL \row2_buffer_reg[164][2]  ( .D(\row2_buffer[165][2] ), .CK(clk), .Q(
        \row2_buffer[164][2] ) );
  DFFQXL \row2_buffer_reg[163][2]  ( .D(\row2_buffer[164][2] ), .CK(clk), .Q(
        \row2_buffer[163][2] ) );
  DFFQXL \row2_buffer_reg[162][2]  ( .D(\row2_buffer[163][2] ), .CK(clk), .Q(
        \row2_buffer[162][2] ) );
  DFFQXL \row2_buffer_reg[161][2]  ( .D(\row2_buffer[162][2] ), .CK(clk), .Q(
        \row2_buffer[161][2] ) );
  DFFQXL \row2_buffer_reg[160][2]  ( .D(\row2_buffer[161][2] ), .CK(clk), .Q(
        \row2_buffer[160][2] ) );
  DFFQXL \row2_buffer_reg[159][2]  ( .D(\row2_buffer[160][2] ), .CK(clk), .Q(
        \row2_buffer[159][2] ) );
  DFFQXL \row2_buffer_reg[158][2]  ( .D(\row2_buffer[159][2] ), .CK(clk), .Q(
        \row2_buffer[158][2] ) );
  DFFQXL \row2_buffer_reg[157][2]  ( .D(\row2_buffer[158][2] ), .CK(clk), .Q(
        \row2_buffer[157][2] ) );
  DFFQXL \row2_buffer_reg[156][2]  ( .D(\row2_buffer[157][2] ), .CK(clk), .Q(
        \row2_buffer[156][2] ) );
  DFFQXL \row2_buffer_reg[155][2]  ( .D(\row2_buffer[156][2] ), .CK(clk), .Q(
        \row2_buffer[155][2] ) );
  DFFQXL \row2_buffer_reg[154][2]  ( .D(\row2_buffer[155][2] ), .CK(clk), .Q(
        \row2_buffer[154][2] ) );
  DFFQXL \row2_buffer_reg[153][2]  ( .D(\row2_buffer[154][2] ), .CK(clk), .Q(
        \row2_buffer[153][2] ) );
  DFFQXL \row2_buffer_reg[152][2]  ( .D(\row2_buffer[153][2] ), .CK(clk), .Q(
        \row2_buffer[152][2] ) );
  DFFQXL \row2_buffer_reg[151][2]  ( .D(\row2_buffer[152][2] ), .CK(clk), .Q(
        \row2_buffer[151][2] ) );
  DFFQXL \row2_buffer_reg[150][2]  ( .D(\row2_buffer[151][2] ), .CK(clk), .Q(
        \row2_buffer[150][2] ) );
  DFFQXL \row2_buffer_reg[149][2]  ( .D(\row2_buffer[150][2] ), .CK(clk), .Q(
        \row2_buffer[149][2] ) );
  DFFQXL \row2_buffer_reg[148][2]  ( .D(\row2_buffer[149][2] ), .CK(clk), .Q(
        \row2_buffer[148][2] ) );
  DFFQXL \row2_buffer_reg[147][2]  ( .D(\row2_buffer[148][2] ), .CK(clk), .Q(
        \row2_buffer[147][2] ) );
  DFFQXL \row2_buffer_reg[146][2]  ( .D(\row2_buffer[147][2] ), .CK(clk), .Q(
        \row2_buffer[146][2] ) );
  DFFQXL \row2_buffer_reg[145][2]  ( .D(\row2_buffer[146][2] ), .CK(clk), .Q(
        \row2_buffer[145][2] ) );
  DFFQXL \row2_buffer_reg[144][2]  ( .D(\row2_buffer[145][2] ), .CK(clk), .Q(
        \row2_buffer[144][2] ) );
  DFFQXL \row2_buffer_reg[143][2]  ( .D(\row2_buffer[144][2] ), .CK(clk), .Q(
        \row2_buffer[143][2] ) );
  DFFQXL \row2_buffer_reg[142][2]  ( .D(\row2_buffer[143][2] ), .CK(clk), .Q(
        \row2_buffer[142][2] ) );
  DFFQXL \row2_buffer_reg[141][2]  ( .D(\row2_buffer[142][2] ), .CK(clk), .Q(
        \row2_buffer[141][2] ) );
  DFFQXL \row2_buffer_reg[140][2]  ( .D(\row2_buffer[141][2] ), .CK(clk), .Q(
        \row2_buffer[140][2] ) );
  DFFQXL \row2_buffer_reg[139][2]  ( .D(\row2_buffer[140][2] ), .CK(clk), .Q(
        \row2_buffer[139][2] ) );
  DFFQXL \row2_buffer_reg[138][2]  ( .D(\row2_buffer[139][2] ), .CK(clk), .Q(
        \row2_buffer[138][2] ) );
  DFFQXL \row2_buffer_reg[137][2]  ( .D(\row2_buffer[138][2] ), .CK(clk), .Q(
        \row2_buffer[137][2] ) );
  DFFQXL \row2_buffer_reg[136][2]  ( .D(\row2_buffer[137][2] ), .CK(clk), .Q(
        \row2_buffer[136][2] ) );
  DFFQXL \row2_buffer_reg[135][2]  ( .D(\row2_buffer[136][2] ), .CK(clk), .Q(
        \row2_buffer[135][2] ) );
  DFFQXL \row2_buffer_reg[134][2]  ( .D(\row2_buffer[135][2] ), .CK(clk), .Q(
        \row2_buffer[134][2] ) );
  DFFQXL \row2_buffer_reg[133][2]  ( .D(\row2_buffer[134][2] ), .CK(clk), .Q(
        \row2_buffer[133][2] ) );
  DFFQXL \row2_buffer_reg[132][2]  ( .D(\row2_buffer[133][2] ), .CK(clk), .Q(
        \row2_buffer[132][2] ) );
  DFFQXL \row2_buffer_reg[131][2]  ( .D(\row2_buffer[132][2] ), .CK(clk), .Q(
        \row2_buffer[131][2] ) );
  DFFQXL \row2_buffer_reg[130][2]  ( .D(\row2_buffer[131][2] ), .CK(clk), .Q(
        \row2_buffer[130][2] ) );
  DFFQXL \row2_buffer_reg[129][2]  ( .D(\row2_buffer[130][2] ), .CK(clk), .Q(
        \row2_buffer[129][2] ) );
  DFFQXL \row2_buffer_reg[128][2]  ( .D(\row2_buffer[129][2] ), .CK(clk), .Q(
        \row2_buffer[128][2] ) );
  DFFQXL \row2_buffer_reg[127][2]  ( .D(\row2_buffer[128][2] ), .CK(clk), .Q(
        \row2_buffer[127][2] ) );
  DFFQXL \row2_buffer_reg[126][2]  ( .D(\row2_buffer[127][2] ), .CK(clk), .Q(
        \row2_buffer[126][2] ) );
  DFFQXL \row2_buffer_reg[125][2]  ( .D(\row2_buffer[126][2] ), .CK(clk), .Q(
        \row2_buffer[125][2] ) );
  DFFQXL \row2_buffer_reg[124][2]  ( .D(\row2_buffer[125][2] ), .CK(clk), .Q(
        \row2_buffer[124][2] ) );
  DFFQXL \row2_buffer_reg[123][2]  ( .D(\row2_buffer[124][2] ), .CK(clk), .Q(
        \row2_buffer[123][2] ) );
  DFFQXL \row2_buffer_reg[122][2]  ( .D(\row2_buffer[123][2] ), .CK(clk), .Q(
        \row2_buffer[122][2] ) );
  DFFQXL \row2_buffer_reg[121][2]  ( .D(\row2_buffer[122][2] ), .CK(clk), .Q(
        \row2_buffer[121][2] ) );
  DFFQXL \row2_buffer_reg[120][2]  ( .D(\row2_buffer[121][2] ), .CK(clk), .Q(
        \row2_buffer[120][2] ) );
  DFFQXL \row2_buffer_reg[119][2]  ( .D(\row2_buffer[120][2] ), .CK(clk), .Q(
        \row2_buffer[119][2] ) );
  DFFQXL \row2_buffer_reg[118][2]  ( .D(\row2_buffer[119][2] ), .CK(clk), .Q(
        \row2_buffer[118][2] ) );
  DFFQXL \row2_buffer_reg[117][2]  ( .D(\row2_buffer[118][2] ), .CK(clk), .Q(
        \row2_buffer[117][2] ) );
  DFFQXL \row2_buffer_reg[116][2]  ( .D(\row2_buffer[117][2] ), .CK(clk), .Q(
        \row2_buffer[116][2] ) );
  DFFQXL \row2_buffer_reg[115][2]  ( .D(\row2_buffer[116][2] ), .CK(clk), .Q(
        \row2_buffer[115][2] ) );
  DFFQXL \row2_buffer_reg[114][2]  ( .D(\row2_buffer[115][2] ), .CK(clk), .Q(
        \row2_buffer[114][2] ) );
  DFFQXL \row2_buffer_reg[113][2]  ( .D(\row2_buffer[114][2] ), .CK(clk), .Q(
        \row2_buffer[113][2] ) );
  DFFQXL \row2_buffer_reg[112][2]  ( .D(\row2_buffer[113][2] ), .CK(clk), .Q(
        \row2_buffer[112][2] ) );
  DFFQXL \row2_buffer_reg[111][2]  ( .D(\row2_buffer[112][2] ), .CK(clk), .Q(
        \row2_buffer[111][2] ) );
  DFFQXL \row2_buffer_reg[110][2]  ( .D(\row2_buffer[111][2] ), .CK(clk), .Q(
        \row2_buffer[110][2] ) );
  DFFQXL \row2_buffer_reg[109][2]  ( .D(\row2_buffer[110][2] ), .CK(clk), .Q(
        \row2_buffer[109][2] ) );
  DFFQXL \row2_buffer_reg[108][2]  ( .D(\row2_buffer[109][2] ), .CK(clk), .Q(
        \row2_buffer[108][2] ) );
  DFFQXL \row2_buffer_reg[107][2]  ( .D(\row2_buffer[108][2] ), .CK(clk), .Q(
        \row2_buffer[107][2] ) );
  DFFQXL \row2_buffer_reg[106][2]  ( .D(\row2_buffer[107][2] ), .CK(clk), .Q(
        \row2_buffer[106][2] ) );
  DFFQXL \row2_buffer_reg[105][2]  ( .D(\row2_buffer[106][2] ), .CK(clk), .Q(
        \row2_buffer[105][2] ) );
  DFFQXL \row2_buffer_reg[104][2]  ( .D(\row2_buffer[105][2] ), .CK(clk), .Q(
        \row2_buffer[104][2] ) );
  DFFQXL \row2_buffer_reg[103][2]  ( .D(\row2_buffer[104][2] ), .CK(clk), .Q(
        \row2_buffer[103][2] ) );
  DFFQXL \row2_buffer_reg[102][2]  ( .D(\row2_buffer[103][2] ), .CK(clk), .Q(
        \row2_buffer[102][2] ) );
  DFFQXL \row2_buffer_reg[101][2]  ( .D(\row2_buffer[102][2] ), .CK(clk), .Q(
        \row2_buffer[101][2] ) );
  DFFQXL \row2_buffer_reg[100][2]  ( .D(\row2_buffer[101][2] ), .CK(clk), .Q(
        \row2_buffer[100][2] ) );
  DFFQXL \row2_buffer_reg[99][2]  ( .D(\row2_buffer[100][2] ), .CK(clk), .Q(
        \row2_buffer[99][2] ) );
  DFFQXL \row2_buffer_reg[98][2]  ( .D(\row2_buffer[99][2] ), .CK(clk), .Q(
        \row2_buffer[98][2] ) );
  DFFQXL \row2_buffer_reg[97][2]  ( .D(\row2_buffer[98][2] ), .CK(clk), .Q(
        \row2_buffer[97][2] ) );
  DFFQXL \row2_buffer_reg[96][2]  ( .D(\row2_buffer[97][2] ), .CK(clk), .Q(
        \row2_buffer[96][2] ) );
  DFFQXL \row2_buffer_reg[95][2]  ( .D(\row2_buffer[96][2] ), .CK(clk), .Q(
        \row2_buffer[95][2] ) );
  DFFQXL \row2_buffer_reg[94][2]  ( .D(\row2_buffer[95][2] ), .CK(clk), .Q(
        \row2_buffer[94][2] ) );
  DFFQXL \row2_buffer_reg[93][2]  ( .D(\row2_buffer[94][2] ), .CK(clk), .Q(
        \row2_buffer[93][2] ) );
  DFFQXL \row2_buffer_reg[92][2]  ( .D(\row2_buffer[93][2] ), .CK(clk), .Q(
        \row2_buffer[92][2] ) );
  DFFQXL \row2_buffer_reg[91][2]  ( .D(\row2_buffer[92][2] ), .CK(clk), .Q(
        \row2_buffer[91][2] ) );
  DFFQXL \row2_buffer_reg[90][2]  ( .D(\row2_buffer[91][2] ), .CK(clk), .Q(
        \row2_buffer[90][2] ) );
  DFFQXL \row2_buffer_reg[89][2]  ( .D(\row2_buffer[90][2] ), .CK(clk), .Q(
        \row2_buffer[89][2] ) );
  DFFQXL \row2_buffer_reg[88][2]  ( .D(\row2_buffer[89][2] ), .CK(clk), .Q(
        \row2_buffer[88][2] ) );
  DFFQXL \row2_buffer_reg[87][2]  ( .D(\row2_buffer[88][2] ), .CK(clk), .Q(
        \row2_buffer[87][2] ) );
  DFFQXL \row2_buffer_reg[86][2]  ( .D(\row2_buffer[87][2] ), .CK(clk), .Q(
        \row2_buffer[86][2] ) );
  DFFQXL \row2_buffer_reg[85][2]  ( .D(\row2_buffer[86][2] ), .CK(clk), .Q(
        \row2_buffer[85][2] ) );
  DFFQXL \row2_buffer_reg[84][2]  ( .D(\row2_buffer[85][2] ), .CK(clk), .Q(
        \row2_buffer[84][2] ) );
  DFFQXL \row2_buffer_reg[83][2]  ( .D(\row2_buffer[84][2] ), .CK(clk), .Q(
        \row2_buffer[83][2] ) );
  DFFQXL \row2_buffer_reg[82][2]  ( .D(\row2_buffer[83][2] ), .CK(clk), .Q(
        \row2_buffer[82][2] ) );
  DFFQXL \row2_buffer_reg[81][2]  ( .D(\row2_buffer[82][2] ), .CK(clk), .Q(
        \row2_buffer[81][2] ) );
  DFFQXL \row2_buffer_reg[80][2]  ( .D(\row2_buffer[81][2] ), .CK(clk), .Q(
        \row2_buffer[80][2] ) );
  DFFQXL \row2_buffer_reg[79][2]  ( .D(\row2_buffer[80][2] ), .CK(clk), .Q(
        \row2_buffer[79][2] ) );
  DFFQXL \row2_buffer_reg[78][2]  ( .D(\row2_buffer[79][2] ), .CK(clk), .Q(
        \row2_buffer[78][2] ) );
  DFFQXL \row2_buffer_reg[77][2]  ( .D(\row2_buffer[78][2] ), .CK(clk), .Q(
        \row2_buffer[77][2] ) );
  DFFQXL \row2_buffer_reg[76][2]  ( .D(\row2_buffer[77][2] ), .CK(clk), .Q(
        \row2_buffer[76][2] ) );
  DFFQXL \row2_buffer_reg[75][2]  ( .D(\row2_buffer[76][2] ), .CK(clk), .Q(
        \row2_buffer[75][2] ) );
  DFFQXL \row2_buffer_reg[74][2]  ( .D(\row2_buffer[75][2] ), .CK(clk), .Q(
        \row2_buffer[74][2] ) );
  DFFQXL \row2_buffer_reg[73][2]  ( .D(\row2_buffer[74][2] ), .CK(clk), .Q(
        \row2_buffer[73][2] ) );
  DFFQXL \row2_buffer_reg[72][2]  ( .D(\row2_buffer[73][2] ), .CK(clk), .Q(
        \row2_buffer[72][2] ) );
  DFFQXL \row2_buffer_reg[71][2]  ( .D(\row2_buffer[72][2] ), .CK(clk), .Q(
        \row2_buffer[71][2] ) );
  DFFQXL \row2_buffer_reg[70][2]  ( .D(\row2_buffer[71][2] ), .CK(clk), .Q(
        \row2_buffer[70][2] ) );
  DFFQXL \row2_buffer_reg[69][2]  ( .D(\row2_buffer[70][2] ), .CK(clk), .Q(
        \row2_buffer[69][2] ) );
  DFFQXL \row2_buffer_reg[68][2]  ( .D(\row2_buffer[69][2] ), .CK(clk), .Q(
        \row2_buffer[68][2] ) );
  DFFQXL \row2_buffer_reg[67][2]  ( .D(\row2_buffer[68][2] ), .CK(clk), .Q(
        \row2_buffer[67][2] ) );
  DFFQXL \row2_buffer_reg[66][2]  ( .D(\row2_buffer[67][2] ), .CK(clk), .Q(
        \row2_buffer[66][2] ) );
  DFFQXL \row2_buffer_reg[65][2]  ( .D(\row2_buffer[66][2] ), .CK(clk), .Q(
        \row2_buffer[65][2] ) );
  DFFQXL \row2_buffer_reg[64][2]  ( .D(\row2_buffer[65][2] ), .CK(clk), .Q(
        \row2_buffer[64][2] ) );
  DFFQXL \row2_buffer_reg[63][2]  ( .D(\row2_buffer[64][2] ), .CK(clk), .Q(
        \row2_buffer[63][2] ) );
  DFFQXL \row2_buffer_reg[62][2]  ( .D(\row2_buffer[63][2] ), .CK(clk), .Q(
        \row2_buffer[62][2] ) );
  DFFQXL \row2_buffer_reg[61][2]  ( .D(\row2_buffer[62][2] ), .CK(clk), .Q(
        \row2_buffer[61][2] ) );
  DFFQXL \row2_buffer_reg[60][2]  ( .D(\row2_buffer[61][2] ), .CK(clk), .Q(
        \row2_buffer[60][2] ) );
  DFFQXL \row2_buffer_reg[59][2]  ( .D(\row2_buffer[60][2] ), .CK(clk), .Q(
        \row2_buffer[59][2] ) );
  DFFQXL \row2_buffer_reg[58][2]  ( .D(\row2_buffer[59][2] ), .CK(clk), .Q(
        \row2_buffer[58][2] ) );
  DFFQXL \row2_buffer_reg[57][2]  ( .D(\row2_buffer[58][2] ), .CK(clk), .Q(
        \row2_buffer[57][2] ) );
  DFFQXL \row2_buffer_reg[56][2]  ( .D(\row2_buffer[57][2] ), .CK(clk), .Q(
        \row2_buffer[56][2] ) );
  DFFQXL \row2_buffer_reg[55][2]  ( .D(\row2_buffer[56][2] ), .CK(clk), .Q(
        \row2_buffer[55][2] ) );
  DFFQXL \row2_buffer_reg[54][2]  ( .D(\row2_buffer[55][2] ), .CK(clk), .Q(
        \row2_buffer[54][2] ) );
  DFFQXL \row2_buffer_reg[53][2]  ( .D(\row2_buffer[54][2] ), .CK(clk), .Q(
        \row2_buffer[53][2] ) );
  DFFQXL \row2_buffer_reg[52][2]  ( .D(\row2_buffer[53][2] ), .CK(clk), .Q(
        \row2_buffer[52][2] ) );
  DFFQXL \row2_buffer_reg[51][2]  ( .D(\row2_buffer[52][2] ), .CK(clk), .Q(
        \row2_buffer[51][2] ) );
  DFFQXL \row2_buffer_reg[50][2]  ( .D(\row2_buffer[51][2] ), .CK(clk), .Q(
        \row2_buffer[50][2] ) );
  DFFQXL \row2_buffer_reg[49][2]  ( .D(\row2_buffer[50][2] ), .CK(clk), .Q(
        \row2_buffer[49][2] ) );
  DFFQXL \row2_buffer_reg[48][2]  ( .D(\row2_buffer[49][2] ), .CK(clk), .Q(
        \row2_buffer[48][2] ) );
  DFFQXL \row2_buffer_reg[47][2]  ( .D(\row2_buffer[48][2] ), .CK(clk), .Q(
        \row2_buffer[47][2] ) );
  DFFQXL \row2_buffer_reg[46][2]  ( .D(\row2_buffer[47][2] ), .CK(clk), .Q(
        \row2_buffer[46][2] ) );
  DFFQXL \row2_buffer_reg[45][2]  ( .D(\row2_buffer[46][2] ), .CK(clk), .Q(
        \row2_buffer[45][2] ) );
  DFFQXL \row2_buffer_reg[44][2]  ( .D(\row2_buffer[45][2] ), .CK(clk), .Q(
        \row2_buffer[44][2] ) );
  DFFQXL \row2_buffer_reg[43][2]  ( .D(\row2_buffer[44][2] ), .CK(clk), .Q(
        \row2_buffer[43][2] ) );
  DFFQXL \row2_buffer_reg[42][2]  ( .D(\row2_buffer[43][2] ), .CK(clk), .Q(
        \row2_buffer[42][2] ) );
  DFFQXL \row2_buffer_reg[41][2]  ( .D(\row2_buffer[42][2] ), .CK(clk), .Q(
        \row2_buffer[41][2] ) );
  DFFQXL \row2_buffer_reg[40][2]  ( .D(\row2_buffer[41][2] ), .CK(clk), .Q(
        \row2_buffer[40][2] ) );
  DFFQXL \row2_buffer_reg[39][2]  ( .D(\row2_buffer[40][2] ), .CK(clk), .Q(
        \row2_buffer[39][2] ) );
  DFFQXL \row2_buffer_reg[38][2]  ( .D(\row2_buffer[39][2] ), .CK(clk), .Q(
        \row2_buffer[38][2] ) );
  DFFQXL \row2_buffer_reg[37][2]  ( .D(\row2_buffer[38][2] ), .CK(clk), .Q(
        \row2_buffer[37][2] ) );
  DFFQXL \row2_buffer_reg[36][2]  ( .D(\row2_buffer[37][2] ), .CK(clk), .Q(
        \row2_buffer[36][2] ) );
  DFFQXL \row2_buffer_reg[35][2]  ( .D(\row2_buffer[36][2] ), .CK(clk), .Q(
        \row2_buffer[35][2] ) );
  DFFQXL \row2_buffer_reg[34][2]  ( .D(\row2_buffer[35][2] ), .CK(clk), .Q(
        \row2_buffer[34][2] ) );
  DFFQXL \row2_buffer_reg[33][2]  ( .D(\row2_buffer[34][2] ), .CK(clk), .Q(
        \row2_buffer[33][2] ) );
  DFFQXL \row2_buffer_reg[32][2]  ( .D(\row2_buffer[33][2] ), .CK(clk), .Q(
        \row2_buffer[32][2] ) );
  DFFQXL \row2_buffer_reg[31][2]  ( .D(\row2_buffer[32][2] ), .CK(clk), .Q(
        \row2_buffer[31][2] ) );
  DFFQXL \row2_buffer_reg[30][2]  ( .D(\row2_buffer[31][2] ), .CK(clk), .Q(
        \row2_buffer[30][2] ) );
  DFFQXL \row2_buffer_reg[29][2]  ( .D(\row2_buffer[30][2] ), .CK(clk), .Q(
        \row2_buffer[29][2] ) );
  DFFQXL \row2_buffer_reg[28][2]  ( .D(\row2_buffer[29][2] ), .CK(clk), .Q(
        \row2_buffer[28][2] ) );
  DFFQXL \row2_buffer_reg[27][2]  ( .D(\row2_buffer[28][2] ), .CK(clk), .Q(
        \row2_buffer[27][2] ) );
  DFFQXL \row2_buffer_reg[26][2]  ( .D(\row2_buffer[27][2] ), .CK(clk), .Q(
        \row2_buffer[26][2] ) );
  DFFQXL \row2_buffer_reg[25][2]  ( .D(\row2_buffer[26][2] ), .CK(clk), .Q(
        \row2_buffer[25][2] ) );
  DFFQXL \row2_buffer_reg[24][2]  ( .D(\row2_buffer[25][2] ), .CK(clk), .Q(
        \row2_buffer[24][2] ) );
  DFFQXL \row2_buffer_reg[23][2]  ( .D(\row2_buffer[24][2] ), .CK(clk), .Q(
        \row2_buffer[23][2] ) );
  DFFQXL \row2_buffer_reg[22][2]  ( .D(\row2_buffer[23][2] ), .CK(clk), .Q(
        \row2_buffer[22][2] ) );
  DFFQXL \row2_buffer_reg[21][2]  ( .D(\row2_buffer[22][2] ), .CK(clk), .Q(
        \row2_buffer[21][2] ) );
  DFFQXL \row2_buffer_reg[20][2]  ( .D(\row2_buffer[21][2] ), .CK(clk), .Q(
        \row2_buffer[20][2] ) );
  DFFQXL \row2_buffer_reg[19][2]  ( .D(\row2_buffer[20][2] ), .CK(clk), .Q(
        \row2_buffer[19][2] ) );
  DFFQXL \row2_buffer_reg[18][2]  ( .D(\row2_buffer[19][2] ), .CK(clk), .Q(
        \row2_buffer[18][2] ) );
  DFFQXL \row2_buffer_reg[17][2]  ( .D(\row2_buffer[18][2] ), .CK(clk), .Q(
        \row2_buffer[17][2] ) );
  DFFQXL \row2_buffer_reg[16][2]  ( .D(\row2_buffer[17][2] ), .CK(clk), .Q(
        \row2_buffer[16][2] ) );
  DFFQXL \row2_buffer_reg[15][2]  ( .D(\row2_buffer[16][2] ), .CK(clk), .Q(
        \row2_buffer[15][2] ) );
  DFFQXL \row2_buffer_reg[14][2]  ( .D(\row2_buffer[15][2] ), .CK(clk), .Q(
        \row2_buffer[14][2] ) );
  DFFQXL \row2_buffer_reg[13][2]  ( .D(\row2_buffer[14][2] ), .CK(clk), .Q(
        \row2_buffer[13][2] ) );
  DFFQXL \row2_buffer_reg[12][2]  ( .D(\row2_buffer[13][2] ), .CK(clk), .Q(
        \row2_buffer[12][2] ) );
  DFFQXL \row2_buffer_reg[11][2]  ( .D(\row2_buffer[12][2] ), .CK(clk), .Q(
        \row2_buffer[11][2] ) );
  DFFQXL \row2_buffer_reg[10][2]  ( .D(\row2_buffer[11][2] ), .CK(clk), .Q(
        \row2_buffer[10][2] ) );
  DFFQXL \row2_buffer_reg[9][2]  ( .D(\row2_buffer[10][2] ), .CK(clk), .Q(
        \row2_buffer[9][2] ) );
  DFFQXL \row2_buffer_reg[8][2]  ( .D(\row2_buffer[9][2] ), .CK(clk), .Q(
        \row2_buffer[8][2] ) );
  DFFQXL \row2_buffer_reg[7][2]  ( .D(\row2_buffer[8][2] ), .CK(clk), .Q(
        \row2_buffer[7][2] ) );
  DFFQXL \row2_buffer_reg[6][2]  ( .D(\row2_buffer[7][2] ), .CK(clk), .Q(
        \row2_buffer[6][2] ) );
  DFFQXL \row2_buffer_reg[5][2]  ( .D(\row2_buffer[6][2] ), .CK(clk), .Q(
        \row2_buffer[5][2] ) );
  DFFQXL \row2_buffer_reg[4][2]  ( .D(\row2_buffer[5][2] ), .CK(clk), .Q(
        \row2_buffer[4][2] ) );
  DFFQXL \row2_buffer_reg[3][2]  ( .D(\row2_buffer[4][2] ), .CK(clk), .Q(
        \row2_buffer[3][2] ) );
  DFFQXL \row1_buffer_reg[225][2]  ( .D(\row2_buffer[0][2] ), .CK(clk), .Q(
        \row1_buffer[225][2] ) );
  DFFQXL \row1_buffer_reg[224][2]  ( .D(\row1_buffer[225][2] ), .CK(clk), .Q(
        \row1_buffer[224][2] ) );
  DFFQXL \row1_buffer_reg[223][2]  ( .D(\row1_buffer[224][2] ), .CK(clk), .Q(
        \row1_buffer[223][2] ) );
  DFFQXL \row1_buffer_reg[222][2]  ( .D(\row1_buffer[223][2] ), .CK(clk), .Q(
        \row1_buffer[222][2] ) );
  DFFQXL \row1_buffer_reg[221][2]  ( .D(\row1_buffer[222][2] ), .CK(clk), .Q(
        \row1_buffer[221][2] ) );
  DFFQXL \row1_buffer_reg[220][2]  ( .D(\row1_buffer[221][2] ), .CK(clk), .Q(
        \row1_buffer[220][2] ) );
  DFFQXL \row1_buffer_reg[219][2]  ( .D(\row1_buffer[220][2] ), .CK(clk), .Q(
        \row1_buffer[219][2] ) );
  DFFQXL \row1_buffer_reg[218][2]  ( .D(\row1_buffer[219][2] ), .CK(clk), .Q(
        \row1_buffer[218][2] ) );
  DFFQXL \row1_buffer_reg[217][2]  ( .D(\row1_buffer[218][2] ), .CK(clk), .Q(
        \row1_buffer[217][2] ) );
  DFFQXL \row1_buffer_reg[216][2]  ( .D(\row1_buffer[217][2] ), .CK(clk), .Q(
        \row1_buffer[216][2] ) );
  DFFQXL \row1_buffer_reg[215][2]  ( .D(\row1_buffer[216][2] ), .CK(clk), .Q(
        \row1_buffer[215][2] ) );
  DFFQXL \row1_buffer_reg[214][2]  ( .D(\row1_buffer[215][2] ), .CK(clk), .Q(
        \row1_buffer[214][2] ) );
  DFFQXL \row1_buffer_reg[213][2]  ( .D(\row1_buffer[214][2] ), .CK(clk), .Q(
        \row1_buffer[213][2] ) );
  DFFQXL \row1_buffer_reg[212][2]  ( .D(\row1_buffer[213][2] ), .CK(clk), .Q(
        \row1_buffer[212][2] ) );
  DFFQXL \row1_buffer_reg[211][2]  ( .D(\row1_buffer[212][2] ), .CK(clk), .Q(
        \row1_buffer[211][2] ) );
  DFFQXL \row1_buffer_reg[210][2]  ( .D(\row1_buffer[211][2] ), .CK(clk), .Q(
        \row1_buffer[210][2] ) );
  DFFQXL \row1_buffer_reg[209][2]  ( .D(\row1_buffer[210][2] ), .CK(clk), .Q(
        \row1_buffer[209][2] ) );
  DFFQXL \row1_buffer_reg[208][2]  ( .D(\row1_buffer[209][2] ), .CK(clk), .Q(
        \row1_buffer[208][2] ) );
  DFFQXL \row1_buffer_reg[207][2]  ( .D(\row1_buffer[208][2] ), .CK(clk), .Q(
        \row1_buffer[207][2] ) );
  DFFQXL \row1_buffer_reg[206][2]  ( .D(\row1_buffer[207][2] ), .CK(clk), .Q(
        \row1_buffer[206][2] ) );
  DFFQXL \row1_buffer_reg[205][2]  ( .D(\row1_buffer[206][2] ), .CK(clk), .Q(
        \row1_buffer[205][2] ) );
  DFFQXL \row1_buffer_reg[204][2]  ( .D(\row1_buffer[205][2] ), .CK(clk), .Q(
        \row1_buffer[204][2] ) );
  DFFQXL \row1_buffer_reg[203][2]  ( .D(\row1_buffer[204][2] ), .CK(clk), .Q(
        \row1_buffer[203][2] ) );
  DFFQXL \row1_buffer_reg[202][2]  ( .D(\row1_buffer[203][2] ), .CK(clk), .Q(
        \row1_buffer[202][2] ) );
  DFFQXL \row1_buffer_reg[201][2]  ( .D(\row1_buffer[202][2] ), .CK(clk), .Q(
        \row1_buffer[201][2] ) );
  DFFQXL \row1_buffer_reg[200][2]  ( .D(\row1_buffer[201][2] ), .CK(clk), .Q(
        \row1_buffer[200][2] ) );
  DFFQXL \row1_buffer_reg[199][2]  ( .D(\row1_buffer[200][2] ), .CK(clk), .Q(
        \row1_buffer[199][2] ) );
  DFFQXL \row1_buffer_reg[198][2]  ( .D(\row1_buffer[199][2] ), .CK(clk), .Q(
        \row1_buffer[198][2] ) );
  DFFQXL \row1_buffer_reg[197][2]  ( .D(\row1_buffer[198][2] ), .CK(clk), .Q(
        \row1_buffer[197][2] ) );
  DFFQXL \row1_buffer_reg[196][2]  ( .D(\row1_buffer[197][2] ), .CK(clk), .Q(
        \row1_buffer[196][2] ) );
  DFFQXL \row1_buffer_reg[195][2]  ( .D(\row1_buffer[196][2] ), .CK(clk), .Q(
        \row1_buffer[195][2] ) );
  DFFQXL \row1_buffer_reg[194][2]  ( .D(\row1_buffer[195][2] ), .CK(clk), .Q(
        \row1_buffer[194][2] ) );
  DFFQXL \row1_buffer_reg[193][2]  ( .D(\row1_buffer[194][2] ), .CK(clk), .Q(
        \row1_buffer[193][2] ) );
  DFFQXL \row1_buffer_reg[192][2]  ( .D(\row1_buffer[193][2] ), .CK(clk), .Q(
        \row1_buffer[192][2] ) );
  DFFQXL \row1_buffer_reg[191][2]  ( .D(\row1_buffer[192][2] ), .CK(clk), .Q(
        \row1_buffer[191][2] ) );
  DFFQXL \row1_buffer_reg[190][2]  ( .D(\row1_buffer[191][2] ), .CK(clk), .Q(
        \row1_buffer[190][2] ) );
  DFFQXL \row1_buffer_reg[189][2]  ( .D(\row1_buffer[190][2] ), .CK(clk), .Q(
        \row1_buffer[189][2] ) );
  DFFQXL \row1_buffer_reg[188][2]  ( .D(\row1_buffer[189][2] ), .CK(clk), .Q(
        \row1_buffer[188][2] ) );
  DFFQXL \row1_buffer_reg[187][2]  ( .D(\row1_buffer[188][2] ), .CK(clk), .Q(
        \row1_buffer[187][2] ) );
  DFFQXL \row1_buffer_reg[186][2]  ( .D(\row1_buffer[187][2] ), .CK(clk), .Q(
        \row1_buffer[186][2] ) );
  DFFQXL \row1_buffer_reg[185][2]  ( .D(\row1_buffer[186][2] ), .CK(clk), .Q(
        \row1_buffer[185][2] ) );
  DFFQXL \row1_buffer_reg[184][2]  ( .D(\row1_buffer[185][2] ), .CK(clk), .Q(
        \row1_buffer[184][2] ) );
  DFFQXL \row1_buffer_reg[183][2]  ( .D(\row1_buffer[184][2] ), .CK(clk), .Q(
        \row1_buffer[183][2] ) );
  DFFQXL \row1_buffer_reg[182][2]  ( .D(\row1_buffer[183][2] ), .CK(clk), .Q(
        \row1_buffer[182][2] ) );
  DFFQXL \row1_buffer_reg[181][2]  ( .D(\row1_buffer[182][2] ), .CK(clk), .Q(
        \row1_buffer[181][2] ) );
  DFFQXL \row1_buffer_reg[180][2]  ( .D(\row1_buffer[181][2] ), .CK(clk), .Q(
        \row1_buffer[180][2] ) );
  DFFQXL \row1_buffer_reg[179][2]  ( .D(\row1_buffer[180][2] ), .CK(clk), .Q(
        \row1_buffer[179][2] ) );
  DFFQXL \row1_buffer_reg[178][2]  ( .D(\row1_buffer[179][2] ), .CK(clk), .Q(
        \row1_buffer[178][2] ) );
  DFFQXL \row1_buffer_reg[177][2]  ( .D(\row1_buffer[178][2] ), .CK(clk), .Q(
        \row1_buffer[177][2] ) );
  DFFQXL \row1_buffer_reg[176][2]  ( .D(\row1_buffer[177][2] ), .CK(clk), .Q(
        \row1_buffer[176][2] ) );
  DFFQXL \row1_buffer_reg[175][2]  ( .D(\row1_buffer[176][2] ), .CK(clk), .Q(
        \row1_buffer[175][2] ) );
  DFFQXL \row1_buffer_reg[174][2]  ( .D(\row1_buffer[175][2] ), .CK(clk), .Q(
        \row1_buffer[174][2] ) );
  DFFQXL \row1_buffer_reg[173][2]  ( .D(\row1_buffer[174][2] ), .CK(clk), .Q(
        \row1_buffer[173][2] ) );
  DFFQXL \row1_buffer_reg[172][2]  ( .D(\row1_buffer[173][2] ), .CK(clk), .Q(
        \row1_buffer[172][2] ) );
  DFFQXL \row1_buffer_reg[171][2]  ( .D(\row1_buffer[172][2] ), .CK(clk), .Q(
        \row1_buffer[171][2] ) );
  DFFQXL \row1_buffer_reg[170][2]  ( .D(\row1_buffer[171][2] ), .CK(clk), .Q(
        \row1_buffer[170][2] ) );
  DFFQXL \row1_buffer_reg[169][2]  ( .D(\row1_buffer[170][2] ), .CK(clk), .Q(
        \row1_buffer[169][2] ) );
  DFFQXL \row1_buffer_reg[168][2]  ( .D(\row1_buffer[169][2] ), .CK(clk), .Q(
        \row1_buffer[168][2] ) );
  DFFQXL \row1_buffer_reg[167][2]  ( .D(\row1_buffer[168][2] ), .CK(clk), .Q(
        \row1_buffer[167][2] ) );
  DFFQXL \row1_buffer_reg[166][2]  ( .D(\row1_buffer[167][2] ), .CK(clk), .Q(
        \row1_buffer[166][2] ) );
  DFFQXL \row1_buffer_reg[165][2]  ( .D(\row1_buffer[166][2] ), .CK(clk), .Q(
        \row1_buffer[165][2] ) );
  DFFQXL \row1_buffer_reg[164][2]  ( .D(\row1_buffer[165][2] ), .CK(clk), .Q(
        \row1_buffer[164][2] ) );
  DFFQXL \row1_buffer_reg[163][2]  ( .D(\row1_buffer[164][2] ), .CK(clk), .Q(
        \row1_buffer[163][2] ) );
  DFFQXL \row1_buffer_reg[162][2]  ( .D(\row1_buffer[163][2] ), .CK(clk), .Q(
        \row1_buffer[162][2] ) );
  DFFQXL \row1_buffer_reg[161][2]  ( .D(\row1_buffer[162][2] ), .CK(clk), .Q(
        \row1_buffer[161][2] ) );
  DFFQXL \row1_buffer_reg[160][2]  ( .D(\row1_buffer[161][2] ), .CK(clk), .Q(
        \row1_buffer[160][2] ) );
  DFFQXL \row1_buffer_reg[159][2]  ( .D(\row1_buffer[160][2] ), .CK(clk), .Q(
        \row1_buffer[159][2] ) );
  DFFQXL \row1_buffer_reg[158][2]  ( .D(\row1_buffer[159][2] ), .CK(clk), .Q(
        \row1_buffer[158][2] ) );
  DFFQXL \row1_buffer_reg[157][2]  ( .D(\row1_buffer[158][2] ), .CK(clk), .Q(
        \row1_buffer[157][2] ) );
  DFFQXL \row1_buffer_reg[156][2]  ( .D(\row1_buffer[157][2] ), .CK(clk), .Q(
        \row1_buffer[156][2] ) );
  DFFQXL \row1_buffer_reg[155][2]  ( .D(\row1_buffer[156][2] ), .CK(clk), .Q(
        \row1_buffer[155][2] ) );
  DFFQXL \row1_buffer_reg[154][2]  ( .D(\row1_buffer[155][2] ), .CK(clk), .Q(
        \row1_buffer[154][2] ) );
  DFFQXL \row1_buffer_reg[153][2]  ( .D(\row1_buffer[154][2] ), .CK(clk), .Q(
        \row1_buffer[153][2] ) );
  DFFQXL \row1_buffer_reg[152][2]  ( .D(\row1_buffer[153][2] ), .CK(clk), .Q(
        \row1_buffer[152][2] ) );
  DFFQXL \row1_buffer_reg[151][2]  ( .D(\row1_buffer[152][2] ), .CK(clk), .Q(
        \row1_buffer[151][2] ) );
  DFFQXL \row1_buffer_reg[150][2]  ( .D(\row1_buffer[151][2] ), .CK(clk), .Q(
        \row1_buffer[150][2] ) );
  DFFQXL \row1_buffer_reg[149][2]  ( .D(\row1_buffer[150][2] ), .CK(clk), .Q(
        \row1_buffer[149][2] ) );
  DFFQXL \row1_buffer_reg[148][2]  ( .D(\row1_buffer[149][2] ), .CK(clk), .Q(
        \row1_buffer[148][2] ) );
  DFFQXL \row1_buffer_reg[147][2]  ( .D(\row1_buffer[148][2] ), .CK(clk), .Q(
        \row1_buffer[147][2] ) );
  DFFQXL \row1_buffer_reg[146][2]  ( .D(\row1_buffer[147][2] ), .CK(clk), .Q(
        \row1_buffer[146][2] ) );
  DFFQXL \row1_buffer_reg[145][2]  ( .D(\row1_buffer[146][2] ), .CK(clk), .Q(
        \row1_buffer[145][2] ) );
  DFFQXL \row1_buffer_reg[144][2]  ( .D(\row1_buffer[145][2] ), .CK(clk), .Q(
        \row1_buffer[144][2] ) );
  DFFQXL \row1_buffer_reg[143][2]  ( .D(\row1_buffer[144][2] ), .CK(clk), .Q(
        \row1_buffer[143][2] ) );
  DFFQXL \row1_buffer_reg[142][2]  ( .D(\row1_buffer[143][2] ), .CK(clk), .Q(
        \row1_buffer[142][2] ) );
  DFFQXL \row1_buffer_reg[141][2]  ( .D(\row1_buffer[142][2] ), .CK(clk), .Q(
        \row1_buffer[141][2] ) );
  DFFQXL \row1_buffer_reg[140][2]  ( .D(\row1_buffer[141][2] ), .CK(clk), .Q(
        \row1_buffer[140][2] ) );
  DFFQXL \row1_buffer_reg[139][2]  ( .D(\row1_buffer[140][2] ), .CK(clk), .Q(
        \row1_buffer[139][2] ) );
  DFFQXL \row1_buffer_reg[138][2]  ( .D(\row1_buffer[139][2] ), .CK(clk), .Q(
        \row1_buffer[138][2] ) );
  DFFQXL \row1_buffer_reg[137][2]  ( .D(\row1_buffer[138][2] ), .CK(clk), .Q(
        \row1_buffer[137][2] ) );
  DFFQXL \row1_buffer_reg[136][2]  ( .D(\row1_buffer[137][2] ), .CK(clk), .Q(
        \row1_buffer[136][2] ) );
  DFFQXL \row1_buffer_reg[135][2]  ( .D(\row1_buffer[136][2] ), .CK(clk), .Q(
        \row1_buffer[135][2] ) );
  DFFQXL \row1_buffer_reg[134][2]  ( .D(\row1_buffer[135][2] ), .CK(clk), .Q(
        \row1_buffer[134][2] ) );
  DFFQXL \row1_buffer_reg[133][2]  ( .D(\row1_buffer[134][2] ), .CK(clk), .Q(
        \row1_buffer[133][2] ) );
  DFFQXL \row1_buffer_reg[132][2]  ( .D(\row1_buffer[133][2] ), .CK(clk), .Q(
        \row1_buffer[132][2] ) );
  DFFQXL \row1_buffer_reg[131][2]  ( .D(\row1_buffer[132][2] ), .CK(clk), .Q(
        \row1_buffer[131][2] ) );
  DFFQXL \row1_buffer_reg[130][2]  ( .D(\row1_buffer[131][2] ), .CK(clk), .Q(
        \row1_buffer[130][2] ) );
  DFFQXL \row1_buffer_reg[129][2]  ( .D(\row1_buffer[130][2] ), .CK(clk), .Q(
        \row1_buffer[129][2] ) );
  DFFQXL \row1_buffer_reg[128][2]  ( .D(\row1_buffer[129][2] ), .CK(clk), .Q(
        \row1_buffer[128][2] ) );
  DFFQXL \row1_buffer_reg[127][2]  ( .D(\row1_buffer[128][2] ), .CK(clk), .Q(
        \row1_buffer[127][2] ) );
  DFFQXL \row1_buffer_reg[126][2]  ( .D(\row1_buffer[127][2] ), .CK(clk), .Q(
        \row1_buffer[126][2] ) );
  DFFQXL \row1_buffer_reg[125][2]  ( .D(\row1_buffer[126][2] ), .CK(clk), .Q(
        \row1_buffer[125][2] ) );
  DFFQXL \row1_buffer_reg[124][2]  ( .D(\row1_buffer[125][2] ), .CK(clk), .Q(
        \row1_buffer[124][2] ) );
  DFFQXL \row1_buffer_reg[123][2]  ( .D(\row1_buffer[124][2] ), .CK(clk), .Q(
        \row1_buffer[123][2] ) );
  DFFQXL \row1_buffer_reg[122][2]  ( .D(\row1_buffer[123][2] ), .CK(clk), .Q(
        \row1_buffer[122][2] ) );
  DFFQXL \row1_buffer_reg[121][2]  ( .D(\row1_buffer[122][2] ), .CK(clk), .Q(
        \row1_buffer[121][2] ) );
  DFFQXL \row1_buffer_reg[120][2]  ( .D(\row1_buffer[121][2] ), .CK(clk), .Q(
        \row1_buffer[120][2] ) );
  DFFQXL \row1_buffer_reg[119][2]  ( .D(\row1_buffer[120][2] ), .CK(clk), .Q(
        \row1_buffer[119][2] ) );
  DFFQXL \row1_buffer_reg[118][2]  ( .D(\row1_buffer[119][2] ), .CK(clk), .Q(
        \row1_buffer[118][2] ) );
  DFFQXL \row1_buffer_reg[117][2]  ( .D(\row1_buffer[118][2] ), .CK(clk), .Q(
        \row1_buffer[117][2] ) );
  DFFQXL \row1_buffer_reg[116][2]  ( .D(\row1_buffer[117][2] ), .CK(clk), .Q(
        \row1_buffer[116][2] ) );
  DFFQXL \row1_buffer_reg[115][2]  ( .D(\row1_buffer[116][2] ), .CK(clk), .Q(
        \row1_buffer[115][2] ) );
  DFFQXL \row1_buffer_reg[114][2]  ( .D(\row1_buffer[115][2] ), .CK(clk), .Q(
        \row1_buffer[114][2] ) );
  DFFQXL \row1_buffer_reg[113][2]  ( .D(\row1_buffer[114][2] ), .CK(clk), .Q(
        \row1_buffer[113][2] ) );
  DFFQXL \row1_buffer_reg[112][2]  ( .D(\row1_buffer[113][2] ), .CK(clk), .Q(
        \row1_buffer[112][2] ) );
  DFFQXL \row1_buffer_reg[111][2]  ( .D(\row1_buffer[112][2] ), .CK(clk), .Q(
        \row1_buffer[111][2] ) );
  DFFQXL \row1_buffer_reg[110][2]  ( .D(\row1_buffer[111][2] ), .CK(clk), .Q(
        \row1_buffer[110][2] ) );
  DFFQXL \row1_buffer_reg[109][2]  ( .D(\row1_buffer[110][2] ), .CK(clk), .Q(
        \row1_buffer[109][2] ) );
  DFFQXL \row1_buffer_reg[108][2]  ( .D(\row1_buffer[109][2] ), .CK(clk), .Q(
        \row1_buffer[108][2] ) );
  DFFQXL \row1_buffer_reg[107][2]  ( .D(\row1_buffer[108][2] ), .CK(clk), .Q(
        \row1_buffer[107][2] ) );
  DFFQXL \row1_buffer_reg[106][2]  ( .D(\row1_buffer[107][2] ), .CK(clk), .Q(
        \row1_buffer[106][2] ) );
  DFFQXL \row1_buffer_reg[105][2]  ( .D(\row1_buffer[106][2] ), .CK(clk), .Q(
        \row1_buffer[105][2] ) );
  DFFQXL \row1_buffer_reg[104][2]  ( .D(\row1_buffer[105][2] ), .CK(clk), .Q(
        \row1_buffer[104][2] ) );
  DFFQXL \row1_buffer_reg[103][2]  ( .D(\row1_buffer[104][2] ), .CK(clk), .Q(
        \row1_buffer[103][2] ) );
  DFFQXL \row1_buffer_reg[102][2]  ( .D(\row1_buffer[103][2] ), .CK(clk), .Q(
        \row1_buffer[102][2] ) );
  DFFQXL \row1_buffer_reg[101][2]  ( .D(\row1_buffer[102][2] ), .CK(clk), .Q(
        \row1_buffer[101][2] ) );
  DFFQXL \row1_buffer_reg[100][2]  ( .D(\row1_buffer[101][2] ), .CK(clk), .Q(
        \row1_buffer[100][2] ) );
  DFFQXL \row1_buffer_reg[99][2]  ( .D(\row1_buffer[100][2] ), .CK(clk), .Q(
        \row1_buffer[99][2] ) );
  DFFQXL \row1_buffer_reg[98][2]  ( .D(\row1_buffer[99][2] ), .CK(clk), .Q(
        \row1_buffer[98][2] ) );
  DFFQXL \row1_buffer_reg[97][2]  ( .D(\row1_buffer[98][2] ), .CK(clk), .Q(
        \row1_buffer[97][2] ) );
  DFFQXL \row1_buffer_reg[96][2]  ( .D(\row1_buffer[97][2] ), .CK(clk), .Q(
        \row1_buffer[96][2] ) );
  DFFQXL \row1_buffer_reg[95][2]  ( .D(\row1_buffer[96][2] ), .CK(clk), .Q(
        \row1_buffer[95][2] ) );
  DFFQXL \row1_buffer_reg[94][2]  ( .D(\row1_buffer[95][2] ), .CK(clk), .Q(
        \row1_buffer[94][2] ) );
  DFFQXL \row1_buffer_reg[93][2]  ( .D(\row1_buffer[94][2] ), .CK(clk), .Q(
        \row1_buffer[93][2] ) );
  DFFQXL \row1_buffer_reg[92][2]  ( .D(\row1_buffer[93][2] ), .CK(clk), .Q(
        \row1_buffer[92][2] ) );
  DFFQXL \row1_buffer_reg[91][2]  ( .D(\row1_buffer[92][2] ), .CK(clk), .Q(
        \row1_buffer[91][2] ) );
  DFFQXL \row1_buffer_reg[90][2]  ( .D(\row1_buffer[91][2] ), .CK(clk), .Q(
        \row1_buffer[90][2] ) );
  DFFQXL \row1_buffer_reg[89][2]  ( .D(\row1_buffer[90][2] ), .CK(clk), .Q(
        \row1_buffer[89][2] ) );
  DFFQXL \row1_buffer_reg[88][2]  ( .D(\row1_buffer[89][2] ), .CK(clk), .Q(
        \row1_buffer[88][2] ) );
  DFFQXL \row1_buffer_reg[87][2]  ( .D(\row1_buffer[88][2] ), .CK(clk), .Q(
        \row1_buffer[87][2] ) );
  DFFQXL \row1_buffer_reg[86][2]  ( .D(\row1_buffer[87][2] ), .CK(clk), .Q(
        \row1_buffer[86][2] ) );
  DFFQXL \row1_buffer_reg[85][2]  ( .D(\row1_buffer[86][2] ), .CK(clk), .Q(
        \row1_buffer[85][2] ) );
  DFFQXL \row1_buffer_reg[84][2]  ( .D(\row1_buffer[85][2] ), .CK(clk), .Q(
        \row1_buffer[84][2] ) );
  DFFQXL \row1_buffer_reg[83][2]  ( .D(\row1_buffer[84][2] ), .CK(clk), .Q(
        \row1_buffer[83][2] ) );
  DFFQXL \row1_buffer_reg[82][2]  ( .D(\row1_buffer[83][2] ), .CK(clk), .Q(
        \row1_buffer[82][2] ) );
  DFFQXL \row1_buffer_reg[81][2]  ( .D(\row1_buffer[82][2] ), .CK(clk), .Q(
        \row1_buffer[81][2] ) );
  DFFQXL \row1_buffer_reg[80][2]  ( .D(\row1_buffer[81][2] ), .CK(clk), .Q(
        \row1_buffer[80][2] ) );
  DFFQXL \row1_buffer_reg[79][2]  ( .D(\row1_buffer[80][2] ), .CK(clk), .Q(
        \row1_buffer[79][2] ) );
  DFFQXL \row1_buffer_reg[78][2]  ( .D(\row1_buffer[79][2] ), .CK(clk), .Q(
        \row1_buffer[78][2] ) );
  DFFQXL \row1_buffer_reg[77][2]  ( .D(\row1_buffer[78][2] ), .CK(clk), .Q(
        \row1_buffer[77][2] ) );
  DFFQXL \row1_buffer_reg[76][2]  ( .D(\row1_buffer[77][2] ), .CK(clk), .Q(
        \row1_buffer[76][2] ) );
  DFFQXL \row1_buffer_reg[75][2]  ( .D(\row1_buffer[76][2] ), .CK(clk), .Q(
        \row1_buffer[75][2] ) );
  DFFQXL \row1_buffer_reg[74][2]  ( .D(\row1_buffer[75][2] ), .CK(clk), .Q(
        \row1_buffer[74][2] ) );
  DFFQXL \row1_buffer_reg[73][2]  ( .D(\row1_buffer[74][2] ), .CK(clk), .Q(
        \row1_buffer[73][2] ) );
  DFFQXL \row1_buffer_reg[72][2]  ( .D(\row1_buffer[73][2] ), .CK(clk), .Q(
        \row1_buffer[72][2] ) );
  DFFQXL \row1_buffer_reg[71][2]  ( .D(\row1_buffer[72][2] ), .CK(clk), .Q(
        \row1_buffer[71][2] ) );
  DFFQXL \row1_buffer_reg[70][2]  ( .D(\row1_buffer[71][2] ), .CK(clk), .Q(
        \row1_buffer[70][2] ) );
  DFFQXL \row1_buffer_reg[69][2]  ( .D(\row1_buffer[70][2] ), .CK(clk), .Q(
        \row1_buffer[69][2] ) );
  DFFQXL \row1_buffer_reg[68][2]  ( .D(\row1_buffer[69][2] ), .CK(clk), .Q(
        \row1_buffer[68][2] ) );
  DFFQXL \row1_buffer_reg[67][2]  ( .D(\row1_buffer[68][2] ), .CK(clk), .Q(
        \row1_buffer[67][2] ) );
  DFFQXL \row1_buffer_reg[66][2]  ( .D(\row1_buffer[67][2] ), .CK(clk), .Q(
        \row1_buffer[66][2] ) );
  DFFQXL \row1_buffer_reg[65][2]  ( .D(\row1_buffer[66][2] ), .CK(clk), .Q(
        \row1_buffer[65][2] ) );
  DFFQXL \row1_buffer_reg[64][2]  ( .D(\row1_buffer[65][2] ), .CK(clk), .Q(
        \row1_buffer[64][2] ) );
  DFFQXL \row1_buffer_reg[63][2]  ( .D(\row1_buffer[64][2] ), .CK(clk), .Q(
        \row1_buffer[63][2] ) );
  DFFQXL \row1_buffer_reg[62][2]  ( .D(\row1_buffer[63][2] ), .CK(clk), .Q(
        \row1_buffer[62][2] ) );
  DFFQXL \row1_buffer_reg[61][2]  ( .D(\row1_buffer[62][2] ), .CK(clk), .Q(
        \row1_buffer[61][2] ) );
  DFFQXL \row1_buffer_reg[60][2]  ( .D(\row1_buffer[61][2] ), .CK(clk), .Q(
        \row1_buffer[60][2] ) );
  DFFQXL \row1_buffer_reg[59][2]  ( .D(\row1_buffer[60][2] ), .CK(clk), .Q(
        \row1_buffer[59][2] ) );
  DFFQXL \row1_buffer_reg[58][2]  ( .D(\row1_buffer[59][2] ), .CK(clk), .Q(
        \row1_buffer[58][2] ) );
  DFFQXL \row1_buffer_reg[57][2]  ( .D(\row1_buffer[58][2] ), .CK(clk), .Q(
        \row1_buffer[57][2] ) );
  DFFQXL \row1_buffer_reg[56][2]  ( .D(\row1_buffer[57][2] ), .CK(clk), .Q(
        \row1_buffer[56][2] ) );
  DFFQXL \row1_buffer_reg[55][2]  ( .D(\row1_buffer[56][2] ), .CK(clk), .Q(
        \row1_buffer[55][2] ) );
  DFFQXL \row1_buffer_reg[54][2]  ( .D(\row1_buffer[55][2] ), .CK(clk), .Q(
        \row1_buffer[54][2] ) );
  DFFQXL \row1_buffer_reg[53][2]  ( .D(\row1_buffer[54][2] ), .CK(clk), .Q(
        \row1_buffer[53][2] ) );
  DFFQXL \row1_buffer_reg[52][2]  ( .D(\row1_buffer[53][2] ), .CK(clk), .Q(
        \row1_buffer[52][2] ) );
  DFFQXL \row1_buffer_reg[51][2]  ( .D(\row1_buffer[52][2] ), .CK(clk), .Q(
        \row1_buffer[51][2] ) );
  DFFQXL \row1_buffer_reg[50][2]  ( .D(\row1_buffer[51][2] ), .CK(clk), .Q(
        \row1_buffer[50][2] ) );
  DFFQXL \row1_buffer_reg[49][2]  ( .D(\row1_buffer[50][2] ), .CK(clk), .Q(
        \row1_buffer[49][2] ) );
  DFFQXL \row1_buffer_reg[48][2]  ( .D(\row1_buffer[49][2] ), .CK(clk), .Q(
        \row1_buffer[48][2] ) );
  DFFQXL \row1_buffer_reg[47][2]  ( .D(\row1_buffer[48][2] ), .CK(clk), .Q(
        \row1_buffer[47][2] ) );
  DFFQXL \row1_buffer_reg[46][2]  ( .D(\row1_buffer[47][2] ), .CK(clk), .Q(
        \row1_buffer[46][2] ) );
  DFFQXL \row1_buffer_reg[45][2]  ( .D(\row1_buffer[46][2] ), .CK(clk), .Q(
        \row1_buffer[45][2] ) );
  DFFQXL \row1_buffer_reg[44][2]  ( .D(\row1_buffer[45][2] ), .CK(clk), .Q(
        \row1_buffer[44][2] ) );
  DFFQXL \row1_buffer_reg[43][2]  ( .D(\row1_buffer[44][2] ), .CK(clk), .Q(
        \row1_buffer[43][2] ) );
  DFFQXL \row1_buffer_reg[42][2]  ( .D(\row1_buffer[43][2] ), .CK(clk), .Q(
        \row1_buffer[42][2] ) );
  DFFQXL \row1_buffer_reg[41][2]  ( .D(\row1_buffer[42][2] ), .CK(clk), .Q(
        \row1_buffer[41][2] ) );
  DFFQXL \row1_buffer_reg[40][2]  ( .D(\row1_buffer[41][2] ), .CK(clk), .Q(
        \row1_buffer[40][2] ) );
  DFFQXL \row1_buffer_reg[39][2]  ( .D(\row1_buffer[40][2] ), .CK(clk), .Q(
        \row1_buffer[39][2] ) );
  DFFQXL \row1_buffer_reg[38][2]  ( .D(\row1_buffer[39][2] ), .CK(clk), .Q(
        \row1_buffer[38][2] ) );
  DFFQXL \row1_buffer_reg[37][2]  ( .D(\row1_buffer[38][2] ), .CK(clk), .Q(
        \row1_buffer[37][2] ) );
  DFFQXL \row1_buffer_reg[36][2]  ( .D(\row1_buffer[37][2] ), .CK(clk), .Q(
        \row1_buffer[36][2] ) );
  DFFQXL \row1_buffer_reg[35][2]  ( .D(\row1_buffer[36][2] ), .CK(clk), .Q(
        \row1_buffer[35][2] ) );
  DFFQXL \row1_buffer_reg[34][2]  ( .D(\row1_buffer[35][2] ), .CK(clk), .Q(
        \row1_buffer[34][2] ) );
  DFFQXL \row1_buffer_reg[33][2]  ( .D(\row1_buffer[34][2] ), .CK(clk), .Q(
        \row1_buffer[33][2] ) );
  DFFQXL \row1_buffer_reg[32][2]  ( .D(\row1_buffer[33][2] ), .CK(clk), .Q(
        \row1_buffer[32][2] ) );
  DFFQXL \row1_buffer_reg[31][2]  ( .D(\row1_buffer[32][2] ), .CK(clk), .Q(
        \row1_buffer[31][2] ) );
  DFFQXL \row1_buffer_reg[30][2]  ( .D(\row1_buffer[31][2] ), .CK(clk), .Q(
        \row1_buffer[30][2] ) );
  DFFQXL \row1_buffer_reg[29][2]  ( .D(\row1_buffer[30][2] ), .CK(clk), .Q(
        \row1_buffer[29][2] ) );
  DFFQXL \row1_buffer_reg[28][2]  ( .D(\row1_buffer[29][2] ), .CK(clk), .Q(
        \row1_buffer[28][2] ) );
  DFFQXL \row1_buffer_reg[27][2]  ( .D(\row1_buffer[28][2] ), .CK(clk), .Q(
        \row1_buffer[27][2] ) );
  DFFQXL \row1_buffer_reg[26][2]  ( .D(\row1_buffer[27][2] ), .CK(clk), .Q(
        \row1_buffer[26][2] ) );
  DFFQXL \row1_buffer_reg[25][2]  ( .D(\row1_buffer[26][2] ), .CK(clk), .Q(
        \row1_buffer[25][2] ) );
  DFFQXL \row1_buffer_reg[24][2]  ( .D(\row1_buffer[25][2] ), .CK(clk), .Q(
        \row1_buffer[24][2] ) );
  DFFQXL \row1_buffer_reg[23][2]  ( .D(\row1_buffer[24][2] ), .CK(clk), .Q(
        \row1_buffer[23][2] ) );
  DFFQXL \row1_buffer_reg[22][2]  ( .D(\row1_buffer[23][2] ), .CK(clk), .Q(
        \row1_buffer[22][2] ) );
  DFFQXL \row1_buffer_reg[21][2]  ( .D(\row1_buffer[22][2] ), .CK(clk), .Q(
        \row1_buffer[21][2] ) );
  DFFQXL \row1_buffer_reg[20][2]  ( .D(\row1_buffer[21][2] ), .CK(clk), .Q(
        \row1_buffer[20][2] ) );
  DFFQXL \row1_buffer_reg[19][2]  ( .D(\row1_buffer[20][2] ), .CK(clk), .Q(
        \row1_buffer[19][2] ) );
  DFFQXL \row1_buffer_reg[18][2]  ( .D(\row1_buffer[19][2] ), .CK(clk), .Q(
        \row1_buffer[18][2] ) );
  DFFQXL \row1_buffer_reg[17][2]  ( .D(\row1_buffer[18][2] ), .CK(clk), .Q(
        \row1_buffer[17][2] ) );
  DFFQXL \row1_buffer_reg[16][2]  ( .D(\row1_buffer[17][2] ), .CK(clk), .Q(
        \row1_buffer[16][2] ) );
  DFFQXL \row1_buffer_reg[15][2]  ( .D(\row1_buffer[16][2] ), .CK(clk), .Q(
        \row1_buffer[15][2] ) );
  DFFQXL \row1_buffer_reg[14][2]  ( .D(\row1_buffer[15][2] ), .CK(clk), .Q(
        \row1_buffer[14][2] ) );
  DFFQXL \row1_buffer_reg[13][2]  ( .D(\row1_buffer[14][2] ), .CK(clk), .Q(
        \row1_buffer[13][2] ) );
  DFFQXL \row1_buffer_reg[12][2]  ( .D(\row1_buffer[13][2] ), .CK(clk), .Q(
        \row1_buffer[12][2] ) );
  DFFQXL \row1_buffer_reg[11][2]  ( .D(\row1_buffer[12][2] ), .CK(clk), .Q(
        \row1_buffer[11][2] ) );
  DFFQXL \row1_buffer_reg[10][2]  ( .D(\row1_buffer[11][2] ), .CK(clk), .Q(
        \row1_buffer[10][2] ) );
  DFFQXL \row1_buffer_reg[9][2]  ( .D(\row1_buffer[10][2] ), .CK(clk), .Q(
        \row1_buffer[9][2] ) );
  DFFQXL \row1_buffer_reg[8][2]  ( .D(\row1_buffer[9][2] ), .CK(clk), .Q(
        \row1_buffer[8][2] ) );
  DFFQXL \row1_buffer_reg[7][2]  ( .D(\row1_buffer[8][2] ), .CK(clk), .Q(
        \row1_buffer[7][2] ) );
  DFFQXL \row1_buffer_reg[6][2]  ( .D(\row1_buffer[7][2] ), .CK(clk), .Q(
        \row1_buffer[6][2] ) );
  DFFQXL \row1_buffer_reg[5][2]  ( .D(\row1_buffer[6][2] ), .CK(clk), .Q(
        \row1_buffer[5][2] ) );
  DFFQXL \row1_buffer_reg[4][2]  ( .D(\row1_buffer[5][2] ), .CK(clk), .Q(
        \row1_buffer[4][2] ) );
  DFFQXL \row1_buffer_reg[3][2]  ( .D(\row1_buffer[4][2] ), .CK(clk), .Q(
        \row1_buffer[3][2] ) );
  DFFQXL \row2_buffer_reg[225][1]  ( .D(\row3_buffer[0][1] ), .CK(clk), .Q(
        \row2_buffer[225][1] ) );
  DFFQXL \row2_buffer_reg[224][1]  ( .D(\row2_buffer[225][1] ), .CK(clk), .Q(
        \row2_buffer[224][1] ) );
  DFFQXL \row2_buffer_reg[223][1]  ( .D(\row2_buffer[224][1] ), .CK(clk), .Q(
        \row2_buffer[223][1] ) );
  DFFQXL \row2_buffer_reg[222][1]  ( .D(\row2_buffer[223][1] ), .CK(clk), .Q(
        \row2_buffer[222][1] ) );
  DFFQXL \row2_buffer_reg[221][1]  ( .D(\row2_buffer[222][1] ), .CK(clk), .Q(
        \row2_buffer[221][1] ) );
  DFFQXL \row2_buffer_reg[220][1]  ( .D(\row2_buffer[221][1] ), .CK(clk), .Q(
        \row2_buffer[220][1] ) );
  DFFQXL \row2_buffer_reg[219][1]  ( .D(\row2_buffer[220][1] ), .CK(clk), .Q(
        \row2_buffer[219][1] ) );
  DFFQXL \row2_buffer_reg[218][1]  ( .D(\row2_buffer[219][1] ), .CK(clk), .Q(
        \row2_buffer[218][1] ) );
  DFFQXL \row2_buffer_reg[217][1]  ( .D(\row2_buffer[218][1] ), .CK(clk), .Q(
        \row2_buffer[217][1] ) );
  DFFQXL \row2_buffer_reg[216][1]  ( .D(\row2_buffer[217][1] ), .CK(clk), .Q(
        \row2_buffer[216][1] ) );
  DFFQXL \row2_buffer_reg[215][1]  ( .D(\row2_buffer[216][1] ), .CK(clk), .Q(
        \row2_buffer[215][1] ) );
  DFFQXL \row2_buffer_reg[214][1]  ( .D(\row2_buffer[215][1] ), .CK(clk), .Q(
        \row2_buffer[214][1] ) );
  DFFQXL \row2_buffer_reg[213][1]  ( .D(\row2_buffer[214][1] ), .CK(clk), .Q(
        \row2_buffer[213][1] ) );
  DFFQXL \row2_buffer_reg[212][1]  ( .D(\row2_buffer[213][1] ), .CK(clk), .Q(
        \row2_buffer[212][1] ) );
  DFFQXL \row2_buffer_reg[211][1]  ( .D(\row2_buffer[212][1] ), .CK(clk), .Q(
        \row2_buffer[211][1] ) );
  DFFQXL \row2_buffer_reg[210][1]  ( .D(\row2_buffer[211][1] ), .CK(clk), .Q(
        \row2_buffer[210][1] ) );
  DFFQXL \row2_buffer_reg[209][1]  ( .D(\row2_buffer[210][1] ), .CK(clk), .Q(
        \row2_buffer[209][1] ) );
  DFFQXL \row2_buffer_reg[208][1]  ( .D(\row2_buffer[209][1] ), .CK(clk), .Q(
        \row2_buffer[208][1] ) );
  DFFQXL \row2_buffer_reg[207][1]  ( .D(\row2_buffer[208][1] ), .CK(clk), .Q(
        \row2_buffer[207][1] ) );
  DFFQXL \row2_buffer_reg[206][1]  ( .D(\row2_buffer[207][1] ), .CK(clk), .Q(
        \row2_buffer[206][1] ) );
  DFFQXL \row2_buffer_reg[205][1]  ( .D(\row2_buffer[206][1] ), .CK(clk), .Q(
        \row2_buffer[205][1] ) );
  DFFQXL \row2_buffer_reg[204][1]  ( .D(\row2_buffer[205][1] ), .CK(clk), .Q(
        \row2_buffer[204][1] ) );
  DFFQXL \row2_buffer_reg[203][1]  ( .D(\row2_buffer[204][1] ), .CK(clk), .Q(
        \row2_buffer[203][1] ) );
  DFFQXL \row2_buffer_reg[202][1]  ( .D(\row2_buffer[203][1] ), .CK(clk), .Q(
        \row2_buffer[202][1] ) );
  DFFQXL \row2_buffer_reg[201][1]  ( .D(\row2_buffer[202][1] ), .CK(clk), .Q(
        \row2_buffer[201][1] ) );
  DFFQXL \row2_buffer_reg[200][1]  ( .D(\row2_buffer[201][1] ), .CK(clk), .Q(
        \row2_buffer[200][1] ) );
  DFFQXL \row2_buffer_reg[199][1]  ( .D(\row2_buffer[200][1] ), .CK(clk), .Q(
        \row2_buffer[199][1] ) );
  DFFQXL \row2_buffer_reg[198][1]  ( .D(\row2_buffer[199][1] ), .CK(clk), .Q(
        \row2_buffer[198][1] ) );
  DFFQXL \row2_buffer_reg[197][1]  ( .D(\row2_buffer[198][1] ), .CK(clk), .Q(
        \row2_buffer[197][1] ) );
  DFFQXL \row2_buffer_reg[196][1]  ( .D(\row2_buffer[197][1] ), .CK(clk), .Q(
        \row2_buffer[196][1] ) );
  DFFQXL \row2_buffer_reg[195][1]  ( .D(\row2_buffer[196][1] ), .CK(clk), .Q(
        \row2_buffer[195][1] ) );
  DFFQXL \row2_buffer_reg[194][1]  ( .D(\row2_buffer[195][1] ), .CK(clk), .Q(
        \row2_buffer[194][1] ) );
  DFFQXL \row2_buffer_reg[193][1]  ( .D(\row2_buffer[194][1] ), .CK(clk), .Q(
        \row2_buffer[193][1] ) );
  DFFQXL \row2_buffer_reg[192][1]  ( .D(\row2_buffer[193][1] ), .CK(clk), .Q(
        \row2_buffer[192][1] ) );
  DFFQXL \row2_buffer_reg[191][1]  ( .D(\row2_buffer[192][1] ), .CK(clk), .Q(
        \row2_buffer[191][1] ) );
  DFFQXL \row2_buffer_reg[190][1]  ( .D(\row2_buffer[191][1] ), .CK(clk), .Q(
        \row2_buffer[190][1] ) );
  DFFQXL \row2_buffer_reg[189][1]  ( .D(\row2_buffer[190][1] ), .CK(clk), .Q(
        \row2_buffer[189][1] ) );
  DFFQXL \row2_buffer_reg[188][1]  ( .D(\row2_buffer[189][1] ), .CK(clk), .Q(
        \row2_buffer[188][1] ) );
  DFFQXL \row2_buffer_reg[187][1]  ( .D(\row2_buffer[188][1] ), .CK(clk), .Q(
        \row2_buffer[187][1] ) );
  DFFQXL \row2_buffer_reg[186][1]  ( .D(\row2_buffer[187][1] ), .CK(clk), .Q(
        \row2_buffer[186][1] ) );
  DFFQXL \row2_buffer_reg[185][1]  ( .D(\row2_buffer[186][1] ), .CK(clk), .Q(
        \row2_buffer[185][1] ) );
  DFFQXL \row2_buffer_reg[184][1]  ( .D(\row2_buffer[185][1] ), .CK(clk), .Q(
        \row2_buffer[184][1] ) );
  DFFQXL \row2_buffer_reg[183][1]  ( .D(\row2_buffer[184][1] ), .CK(clk), .Q(
        \row2_buffer[183][1] ) );
  DFFQXL \row2_buffer_reg[182][1]  ( .D(\row2_buffer[183][1] ), .CK(clk), .Q(
        \row2_buffer[182][1] ) );
  DFFQXL \row2_buffer_reg[181][1]  ( .D(\row2_buffer[182][1] ), .CK(clk), .Q(
        \row2_buffer[181][1] ) );
  DFFQXL \row2_buffer_reg[180][1]  ( .D(\row2_buffer[181][1] ), .CK(clk), .Q(
        \row2_buffer[180][1] ) );
  DFFQXL \row2_buffer_reg[179][1]  ( .D(\row2_buffer[180][1] ), .CK(clk), .Q(
        \row2_buffer[179][1] ) );
  DFFQXL \row2_buffer_reg[178][1]  ( .D(\row2_buffer[179][1] ), .CK(clk), .Q(
        \row2_buffer[178][1] ) );
  DFFQXL \row2_buffer_reg[177][1]  ( .D(\row2_buffer[178][1] ), .CK(clk), .Q(
        \row2_buffer[177][1] ) );
  DFFQXL \row2_buffer_reg[176][1]  ( .D(\row2_buffer[177][1] ), .CK(clk), .Q(
        \row2_buffer[176][1] ) );
  DFFQXL \row2_buffer_reg[175][1]  ( .D(\row2_buffer[176][1] ), .CK(clk), .Q(
        \row2_buffer[175][1] ) );
  DFFQXL \row2_buffer_reg[174][1]  ( .D(\row2_buffer[175][1] ), .CK(clk), .Q(
        \row2_buffer[174][1] ) );
  DFFQXL \row2_buffer_reg[173][1]  ( .D(\row2_buffer[174][1] ), .CK(clk), .Q(
        \row2_buffer[173][1] ) );
  DFFQXL \row2_buffer_reg[172][1]  ( .D(\row2_buffer[173][1] ), .CK(clk), .Q(
        \row2_buffer[172][1] ) );
  DFFQXL \row2_buffer_reg[171][1]  ( .D(\row2_buffer[172][1] ), .CK(clk), .Q(
        \row2_buffer[171][1] ) );
  DFFQXL \row2_buffer_reg[170][1]  ( .D(\row2_buffer[171][1] ), .CK(clk), .Q(
        \row2_buffer[170][1] ) );
  DFFQXL \row2_buffer_reg[169][1]  ( .D(\row2_buffer[170][1] ), .CK(clk), .Q(
        \row2_buffer[169][1] ) );
  DFFQXL \row2_buffer_reg[168][1]  ( .D(\row2_buffer[169][1] ), .CK(clk), .Q(
        \row2_buffer[168][1] ) );
  DFFQXL \row2_buffer_reg[167][1]  ( .D(\row2_buffer[168][1] ), .CK(clk), .Q(
        \row2_buffer[167][1] ) );
  DFFQXL \row2_buffer_reg[166][1]  ( .D(\row2_buffer[167][1] ), .CK(clk), .Q(
        \row2_buffer[166][1] ) );
  DFFQXL \row2_buffer_reg[165][1]  ( .D(\row2_buffer[166][1] ), .CK(clk), .Q(
        \row2_buffer[165][1] ) );
  DFFQXL \row2_buffer_reg[164][1]  ( .D(\row2_buffer[165][1] ), .CK(clk), .Q(
        \row2_buffer[164][1] ) );
  DFFQXL \row2_buffer_reg[163][1]  ( .D(\row2_buffer[164][1] ), .CK(clk), .Q(
        \row2_buffer[163][1] ) );
  DFFQXL \row2_buffer_reg[162][1]  ( .D(\row2_buffer[163][1] ), .CK(clk), .Q(
        \row2_buffer[162][1] ) );
  DFFQXL \row2_buffer_reg[161][1]  ( .D(\row2_buffer[162][1] ), .CK(clk), .Q(
        \row2_buffer[161][1] ) );
  DFFQXL \row2_buffer_reg[160][1]  ( .D(\row2_buffer[161][1] ), .CK(clk), .Q(
        \row2_buffer[160][1] ) );
  DFFQXL \row2_buffer_reg[159][1]  ( .D(\row2_buffer[160][1] ), .CK(clk), .Q(
        \row2_buffer[159][1] ) );
  DFFQXL \row2_buffer_reg[158][1]  ( .D(\row2_buffer[159][1] ), .CK(clk), .Q(
        \row2_buffer[158][1] ) );
  DFFQXL \row2_buffer_reg[157][1]  ( .D(\row2_buffer[158][1] ), .CK(clk), .Q(
        \row2_buffer[157][1] ) );
  DFFQXL \row2_buffer_reg[156][1]  ( .D(\row2_buffer[157][1] ), .CK(clk), .Q(
        \row2_buffer[156][1] ) );
  DFFQXL \row2_buffer_reg[155][1]  ( .D(\row2_buffer[156][1] ), .CK(clk), .Q(
        \row2_buffer[155][1] ) );
  DFFQXL \row2_buffer_reg[154][1]  ( .D(\row2_buffer[155][1] ), .CK(clk), .Q(
        \row2_buffer[154][1] ) );
  DFFQXL \row2_buffer_reg[153][1]  ( .D(\row2_buffer[154][1] ), .CK(clk), .Q(
        \row2_buffer[153][1] ) );
  DFFQXL \row2_buffer_reg[152][1]  ( .D(\row2_buffer[153][1] ), .CK(clk), .Q(
        \row2_buffer[152][1] ) );
  DFFQXL \row2_buffer_reg[151][1]  ( .D(\row2_buffer[152][1] ), .CK(clk), .Q(
        \row2_buffer[151][1] ) );
  DFFQXL \row2_buffer_reg[150][1]  ( .D(\row2_buffer[151][1] ), .CK(clk), .Q(
        \row2_buffer[150][1] ) );
  DFFQXL \row2_buffer_reg[149][1]  ( .D(\row2_buffer[150][1] ), .CK(clk), .Q(
        \row2_buffer[149][1] ) );
  DFFQXL \row2_buffer_reg[148][1]  ( .D(\row2_buffer[149][1] ), .CK(clk), .Q(
        \row2_buffer[148][1] ) );
  DFFQXL \row2_buffer_reg[147][1]  ( .D(\row2_buffer[148][1] ), .CK(clk), .Q(
        \row2_buffer[147][1] ) );
  DFFQXL \row2_buffer_reg[146][1]  ( .D(\row2_buffer[147][1] ), .CK(clk), .Q(
        \row2_buffer[146][1] ) );
  DFFQXL \row2_buffer_reg[145][1]  ( .D(\row2_buffer[146][1] ), .CK(clk), .Q(
        \row2_buffer[145][1] ) );
  DFFQXL \row2_buffer_reg[144][1]  ( .D(\row2_buffer[145][1] ), .CK(clk), .Q(
        \row2_buffer[144][1] ) );
  DFFQXL \row2_buffer_reg[143][1]  ( .D(\row2_buffer[144][1] ), .CK(clk), .Q(
        \row2_buffer[143][1] ) );
  DFFQXL \row2_buffer_reg[142][1]  ( .D(\row2_buffer[143][1] ), .CK(clk), .Q(
        \row2_buffer[142][1] ) );
  DFFQXL \row2_buffer_reg[141][1]  ( .D(\row2_buffer[142][1] ), .CK(clk), .Q(
        \row2_buffer[141][1] ) );
  DFFQXL \row2_buffer_reg[140][1]  ( .D(\row2_buffer[141][1] ), .CK(clk), .Q(
        \row2_buffer[140][1] ) );
  DFFQXL \row2_buffer_reg[139][1]  ( .D(\row2_buffer[140][1] ), .CK(clk), .Q(
        \row2_buffer[139][1] ) );
  DFFQXL \row2_buffer_reg[138][1]  ( .D(\row2_buffer[139][1] ), .CK(clk), .Q(
        \row2_buffer[138][1] ) );
  DFFQXL \row2_buffer_reg[137][1]  ( .D(\row2_buffer[138][1] ), .CK(clk), .Q(
        \row2_buffer[137][1] ) );
  DFFQXL \row2_buffer_reg[136][1]  ( .D(\row2_buffer[137][1] ), .CK(clk), .Q(
        \row2_buffer[136][1] ) );
  DFFQXL \row2_buffer_reg[135][1]  ( .D(\row2_buffer[136][1] ), .CK(clk), .Q(
        \row2_buffer[135][1] ) );
  DFFQXL \row2_buffer_reg[134][1]  ( .D(\row2_buffer[135][1] ), .CK(clk), .Q(
        \row2_buffer[134][1] ) );
  DFFQXL \row2_buffer_reg[133][1]  ( .D(\row2_buffer[134][1] ), .CK(clk), .Q(
        \row2_buffer[133][1] ) );
  DFFQXL \row2_buffer_reg[132][1]  ( .D(\row2_buffer[133][1] ), .CK(clk), .Q(
        \row2_buffer[132][1] ) );
  DFFQXL \row2_buffer_reg[131][1]  ( .D(\row2_buffer[132][1] ), .CK(clk), .Q(
        \row2_buffer[131][1] ) );
  DFFQXL \row2_buffer_reg[130][1]  ( .D(\row2_buffer[131][1] ), .CK(clk), .Q(
        \row2_buffer[130][1] ) );
  DFFQXL \row2_buffer_reg[129][1]  ( .D(\row2_buffer[130][1] ), .CK(clk), .Q(
        \row2_buffer[129][1] ) );
  DFFQXL \row2_buffer_reg[128][1]  ( .D(\row2_buffer[129][1] ), .CK(clk), .Q(
        \row2_buffer[128][1] ) );
  DFFQXL \row2_buffer_reg[127][1]  ( .D(\row2_buffer[128][1] ), .CK(clk), .Q(
        \row2_buffer[127][1] ) );
  DFFQXL \row2_buffer_reg[126][1]  ( .D(\row2_buffer[127][1] ), .CK(clk), .Q(
        \row2_buffer[126][1] ) );
  DFFQXL \row2_buffer_reg[125][1]  ( .D(\row2_buffer[126][1] ), .CK(clk), .Q(
        \row2_buffer[125][1] ) );
  DFFQXL \row2_buffer_reg[124][1]  ( .D(\row2_buffer[125][1] ), .CK(clk), .Q(
        \row2_buffer[124][1] ) );
  DFFQXL \row2_buffer_reg[123][1]  ( .D(\row2_buffer[124][1] ), .CK(clk), .Q(
        \row2_buffer[123][1] ) );
  DFFQXL \row2_buffer_reg[122][1]  ( .D(\row2_buffer[123][1] ), .CK(clk), .Q(
        \row2_buffer[122][1] ) );
  DFFQXL \row2_buffer_reg[121][1]  ( .D(\row2_buffer[122][1] ), .CK(clk), .Q(
        \row2_buffer[121][1] ) );
  DFFQXL \row2_buffer_reg[120][1]  ( .D(\row2_buffer[121][1] ), .CK(clk), .Q(
        \row2_buffer[120][1] ) );
  DFFQXL \row2_buffer_reg[119][1]  ( .D(\row2_buffer[120][1] ), .CK(clk), .Q(
        \row2_buffer[119][1] ) );
  DFFQXL \row2_buffer_reg[118][1]  ( .D(\row2_buffer[119][1] ), .CK(clk), .Q(
        \row2_buffer[118][1] ) );
  DFFQXL \row2_buffer_reg[117][1]  ( .D(\row2_buffer[118][1] ), .CK(clk), .Q(
        \row2_buffer[117][1] ) );
  DFFQXL \row2_buffer_reg[116][1]  ( .D(\row2_buffer[117][1] ), .CK(clk), .Q(
        \row2_buffer[116][1] ) );
  DFFQXL \row2_buffer_reg[115][1]  ( .D(\row2_buffer[116][1] ), .CK(clk), .Q(
        \row2_buffer[115][1] ) );
  DFFQXL \row2_buffer_reg[114][1]  ( .D(\row2_buffer[115][1] ), .CK(clk), .Q(
        \row2_buffer[114][1] ) );
  DFFQXL \row2_buffer_reg[113][1]  ( .D(\row2_buffer[114][1] ), .CK(clk), .Q(
        \row2_buffer[113][1] ) );
  DFFQXL \row2_buffer_reg[112][1]  ( .D(\row2_buffer[113][1] ), .CK(clk), .Q(
        \row2_buffer[112][1] ) );
  DFFQXL \row2_buffer_reg[111][1]  ( .D(\row2_buffer[112][1] ), .CK(clk), .Q(
        \row2_buffer[111][1] ) );
  DFFQXL \row2_buffer_reg[110][1]  ( .D(\row2_buffer[111][1] ), .CK(clk), .Q(
        \row2_buffer[110][1] ) );
  DFFQXL \row2_buffer_reg[109][1]  ( .D(\row2_buffer[110][1] ), .CK(clk), .Q(
        \row2_buffer[109][1] ) );
  DFFQXL \row2_buffer_reg[108][1]  ( .D(\row2_buffer[109][1] ), .CK(clk), .Q(
        \row2_buffer[108][1] ) );
  DFFQXL \row2_buffer_reg[107][1]  ( .D(\row2_buffer[108][1] ), .CK(clk), .Q(
        \row2_buffer[107][1] ) );
  DFFQXL \row2_buffer_reg[106][1]  ( .D(\row2_buffer[107][1] ), .CK(clk), .Q(
        \row2_buffer[106][1] ) );
  DFFQXL \row2_buffer_reg[105][1]  ( .D(\row2_buffer[106][1] ), .CK(clk), .Q(
        \row2_buffer[105][1] ) );
  DFFQXL \row2_buffer_reg[104][1]  ( .D(\row2_buffer[105][1] ), .CK(clk), .Q(
        \row2_buffer[104][1] ) );
  DFFQXL \row2_buffer_reg[103][1]  ( .D(\row2_buffer[104][1] ), .CK(clk), .Q(
        \row2_buffer[103][1] ) );
  DFFQXL \row2_buffer_reg[102][1]  ( .D(\row2_buffer[103][1] ), .CK(clk), .Q(
        \row2_buffer[102][1] ) );
  DFFQXL \row2_buffer_reg[101][1]  ( .D(\row2_buffer[102][1] ), .CK(clk), .Q(
        \row2_buffer[101][1] ) );
  DFFQXL \row2_buffer_reg[100][1]  ( .D(\row2_buffer[101][1] ), .CK(clk), .Q(
        \row2_buffer[100][1] ) );
  DFFQXL \row2_buffer_reg[99][1]  ( .D(\row2_buffer[100][1] ), .CK(clk), .Q(
        \row2_buffer[99][1] ) );
  DFFQXL \row2_buffer_reg[98][1]  ( .D(\row2_buffer[99][1] ), .CK(clk), .Q(
        \row2_buffer[98][1] ) );
  DFFQXL \row2_buffer_reg[97][1]  ( .D(\row2_buffer[98][1] ), .CK(clk), .Q(
        \row2_buffer[97][1] ) );
  DFFQXL \row2_buffer_reg[96][1]  ( .D(\row2_buffer[97][1] ), .CK(clk), .Q(
        \row2_buffer[96][1] ) );
  DFFQXL \row2_buffer_reg[95][1]  ( .D(\row2_buffer[96][1] ), .CK(clk), .Q(
        \row2_buffer[95][1] ) );
  DFFQXL \row2_buffer_reg[94][1]  ( .D(\row2_buffer[95][1] ), .CK(clk), .Q(
        \row2_buffer[94][1] ) );
  DFFQXL \row2_buffer_reg[93][1]  ( .D(\row2_buffer[94][1] ), .CK(clk), .Q(
        \row2_buffer[93][1] ) );
  DFFQXL \row2_buffer_reg[92][1]  ( .D(\row2_buffer[93][1] ), .CK(clk), .Q(
        \row2_buffer[92][1] ) );
  DFFQXL \row2_buffer_reg[91][1]  ( .D(\row2_buffer[92][1] ), .CK(clk), .Q(
        \row2_buffer[91][1] ) );
  DFFQXL \row2_buffer_reg[90][1]  ( .D(\row2_buffer[91][1] ), .CK(clk), .Q(
        \row2_buffer[90][1] ) );
  DFFQXL \row2_buffer_reg[89][1]  ( .D(\row2_buffer[90][1] ), .CK(clk), .Q(
        \row2_buffer[89][1] ) );
  DFFQXL \row2_buffer_reg[88][1]  ( .D(\row2_buffer[89][1] ), .CK(clk), .Q(
        \row2_buffer[88][1] ) );
  DFFQXL \row2_buffer_reg[87][1]  ( .D(\row2_buffer[88][1] ), .CK(clk), .Q(
        \row2_buffer[87][1] ) );
  DFFQXL \row2_buffer_reg[86][1]  ( .D(\row2_buffer[87][1] ), .CK(clk), .Q(
        \row2_buffer[86][1] ) );
  DFFQXL \row2_buffer_reg[85][1]  ( .D(\row2_buffer[86][1] ), .CK(clk), .Q(
        \row2_buffer[85][1] ) );
  DFFQXL \row2_buffer_reg[84][1]  ( .D(\row2_buffer[85][1] ), .CK(clk), .Q(
        \row2_buffer[84][1] ) );
  DFFQXL \row2_buffer_reg[83][1]  ( .D(\row2_buffer[84][1] ), .CK(clk), .Q(
        \row2_buffer[83][1] ) );
  DFFQXL \row2_buffer_reg[82][1]  ( .D(\row2_buffer[83][1] ), .CK(clk), .Q(
        \row2_buffer[82][1] ) );
  DFFQXL \row2_buffer_reg[81][1]  ( .D(\row2_buffer[82][1] ), .CK(clk), .Q(
        \row2_buffer[81][1] ) );
  DFFQXL \row2_buffer_reg[80][1]  ( .D(\row2_buffer[81][1] ), .CK(clk), .Q(
        \row2_buffer[80][1] ) );
  DFFQXL \row2_buffer_reg[79][1]  ( .D(\row2_buffer[80][1] ), .CK(clk), .Q(
        \row2_buffer[79][1] ) );
  DFFQXL \row2_buffer_reg[78][1]  ( .D(\row2_buffer[79][1] ), .CK(clk), .Q(
        \row2_buffer[78][1] ) );
  DFFQXL \row2_buffer_reg[77][1]  ( .D(\row2_buffer[78][1] ), .CK(clk), .Q(
        \row2_buffer[77][1] ) );
  DFFQXL \row2_buffer_reg[76][1]  ( .D(\row2_buffer[77][1] ), .CK(clk), .Q(
        \row2_buffer[76][1] ) );
  DFFQXL \row2_buffer_reg[75][1]  ( .D(\row2_buffer[76][1] ), .CK(clk), .Q(
        \row2_buffer[75][1] ) );
  DFFQXL \row2_buffer_reg[74][1]  ( .D(\row2_buffer[75][1] ), .CK(clk), .Q(
        \row2_buffer[74][1] ) );
  DFFQXL \row2_buffer_reg[73][1]  ( .D(\row2_buffer[74][1] ), .CK(clk), .Q(
        \row2_buffer[73][1] ) );
  DFFQXL \row2_buffer_reg[72][1]  ( .D(\row2_buffer[73][1] ), .CK(clk), .Q(
        \row2_buffer[72][1] ) );
  DFFQXL \row2_buffer_reg[71][1]  ( .D(\row2_buffer[72][1] ), .CK(clk), .Q(
        \row2_buffer[71][1] ) );
  DFFQXL \row2_buffer_reg[70][1]  ( .D(\row2_buffer[71][1] ), .CK(clk), .Q(
        \row2_buffer[70][1] ) );
  DFFQXL \row2_buffer_reg[69][1]  ( .D(\row2_buffer[70][1] ), .CK(clk), .Q(
        \row2_buffer[69][1] ) );
  DFFQXL \row2_buffer_reg[68][1]  ( .D(\row2_buffer[69][1] ), .CK(clk), .Q(
        \row2_buffer[68][1] ) );
  DFFQXL \row2_buffer_reg[67][1]  ( .D(\row2_buffer[68][1] ), .CK(clk), .Q(
        \row2_buffer[67][1] ) );
  DFFQXL \row2_buffer_reg[66][1]  ( .D(\row2_buffer[67][1] ), .CK(clk), .Q(
        \row2_buffer[66][1] ) );
  DFFQXL \row2_buffer_reg[65][1]  ( .D(\row2_buffer[66][1] ), .CK(clk), .Q(
        \row2_buffer[65][1] ) );
  DFFQXL \row2_buffer_reg[64][1]  ( .D(\row2_buffer[65][1] ), .CK(clk), .Q(
        \row2_buffer[64][1] ) );
  DFFQXL \row2_buffer_reg[63][1]  ( .D(\row2_buffer[64][1] ), .CK(clk), .Q(
        \row2_buffer[63][1] ) );
  DFFQXL \row2_buffer_reg[62][1]  ( .D(\row2_buffer[63][1] ), .CK(clk), .Q(
        \row2_buffer[62][1] ) );
  DFFQXL \row2_buffer_reg[61][1]  ( .D(\row2_buffer[62][1] ), .CK(clk), .Q(
        \row2_buffer[61][1] ) );
  DFFQXL \row2_buffer_reg[60][1]  ( .D(\row2_buffer[61][1] ), .CK(clk), .Q(
        \row2_buffer[60][1] ) );
  DFFQXL \row2_buffer_reg[59][1]  ( .D(\row2_buffer[60][1] ), .CK(clk), .Q(
        \row2_buffer[59][1] ) );
  DFFQXL \row2_buffer_reg[58][1]  ( .D(\row2_buffer[59][1] ), .CK(clk), .Q(
        \row2_buffer[58][1] ) );
  DFFQXL \row2_buffer_reg[57][1]  ( .D(\row2_buffer[58][1] ), .CK(clk), .Q(
        \row2_buffer[57][1] ) );
  DFFQXL \row2_buffer_reg[56][1]  ( .D(\row2_buffer[57][1] ), .CK(clk), .Q(
        \row2_buffer[56][1] ) );
  DFFQXL \row2_buffer_reg[55][1]  ( .D(\row2_buffer[56][1] ), .CK(clk), .Q(
        \row2_buffer[55][1] ) );
  DFFQXL \row2_buffer_reg[54][1]  ( .D(\row2_buffer[55][1] ), .CK(clk), .Q(
        \row2_buffer[54][1] ) );
  DFFQXL \row2_buffer_reg[53][1]  ( .D(\row2_buffer[54][1] ), .CK(clk), .Q(
        \row2_buffer[53][1] ) );
  DFFQXL \row2_buffer_reg[52][1]  ( .D(\row2_buffer[53][1] ), .CK(clk), .Q(
        \row2_buffer[52][1] ) );
  DFFQXL \row2_buffer_reg[51][1]  ( .D(\row2_buffer[52][1] ), .CK(clk), .Q(
        \row2_buffer[51][1] ) );
  DFFQXL \row2_buffer_reg[50][1]  ( .D(\row2_buffer[51][1] ), .CK(clk), .Q(
        \row2_buffer[50][1] ) );
  DFFQXL \row2_buffer_reg[49][1]  ( .D(\row2_buffer[50][1] ), .CK(clk), .Q(
        \row2_buffer[49][1] ) );
  DFFQXL \row2_buffer_reg[48][1]  ( .D(\row2_buffer[49][1] ), .CK(clk), .Q(
        \row2_buffer[48][1] ) );
  DFFQXL \row2_buffer_reg[47][1]  ( .D(\row2_buffer[48][1] ), .CK(clk), .Q(
        \row2_buffer[47][1] ) );
  DFFQXL \row2_buffer_reg[46][1]  ( .D(\row2_buffer[47][1] ), .CK(clk), .Q(
        \row2_buffer[46][1] ) );
  DFFQXL \row2_buffer_reg[45][1]  ( .D(\row2_buffer[46][1] ), .CK(clk), .Q(
        \row2_buffer[45][1] ) );
  DFFQXL \row2_buffer_reg[44][1]  ( .D(\row2_buffer[45][1] ), .CK(clk), .Q(
        \row2_buffer[44][1] ) );
  DFFQXL \row2_buffer_reg[43][1]  ( .D(\row2_buffer[44][1] ), .CK(clk), .Q(
        \row2_buffer[43][1] ) );
  DFFQXL \row2_buffer_reg[42][1]  ( .D(\row2_buffer[43][1] ), .CK(clk), .Q(
        \row2_buffer[42][1] ) );
  DFFQXL \row2_buffer_reg[41][1]  ( .D(\row2_buffer[42][1] ), .CK(clk), .Q(
        \row2_buffer[41][1] ) );
  DFFQXL \row2_buffer_reg[40][1]  ( .D(\row2_buffer[41][1] ), .CK(clk), .Q(
        \row2_buffer[40][1] ) );
  DFFQXL \row2_buffer_reg[39][1]  ( .D(\row2_buffer[40][1] ), .CK(clk), .Q(
        \row2_buffer[39][1] ) );
  DFFQXL \row2_buffer_reg[38][1]  ( .D(\row2_buffer[39][1] ), .CK(clk), .Q(
        \row2_buffer[38][1] ) );
  DFFQXL \row2_buffer_reg[37][1]  ( .D(\row2_buffer[38][1] ), .CK(clk), .Q(
        \row2_buffer[37][1] ) );
  DFFQXL \row2_buffer_reg[36][1]  ( .D(\row2_buffer[37][1] ), .CK(clk), .Q(
        \row2_buffer[36][1] ) );
  DFFQXL \row2_buffer_reg[35][1]  ( .D(\row2_buffer[36][1] ), .CK(clk), .Q(
        \row2_buffer[35][1] ) );
  DFFQXL \row2_buffer_reg[34][1]  ( .D(\row2_buffer[35][1] ), .CK(clk), .Q(
        \row2_buffer[34][1] ) );
  DFFQXL \row2_buffer_reg[33][1]  ( .D(\row2_buffer[34][1] ), .CK(clk), .Q(
        \row2_buffer[33][1] ) );
  DFFQXL \row2_buffer_reg[32][1]  ( .D(\row2_buffer[33][1] ), .CK(clk), .Q(
        \row2_buffer[32][1] ) );
  DFFQXL \row2_buffer_reg[31][1]  ( .D(\row2_buffer[32][1] ), .CK(clk), .Q(
        \row2_buffer[31][1] ) );
  DFFQXL \row2_buffer_reg[30][1]  ( .D(\row2_buffer[31][1] ), .CK(clk), .Q(
        \row2_buffer[30][1] ) );
  DFFQXL \row2_buffer_reg[29][1]  ( .D(\row2_buffer[30][1] ), .CK(clk), .Q(
        \row2_buffer[29][1] ) );
  DFFQXL \row2_buffer_reg[28][1]  ( .D(\row2_buffer[29][1] ), .CK(clk), .Q(
        \row2_buffer[28][1] ) );
  DFFQXL \row2_buffer_reg[27][1]  ( .D(\row2_buffer[28][1] ), .CK(clk), .Q(
        \row2_buffer[27][1] ) );
  DFFQXL \row2_buffer_reg[26][1]  ( .D(\row2_buffer[27][1] ), .CK(clk), .Q(
        \row2_buffer[26][1] ) );
  DFFQXL \row2_buffer_reg[25][1]  ( .D(\row2_buffer[26][1] ), .CK(clk), .Q(
        \row2_buffer[25][1] ) );
  DFFQXL \row2_buffer_reg[24][1]  ( .D(\row2_buffer[25][1] ), .CK(clk), .Q(
        \row2_buffer[24][1] ) );
  DFFQXL \row2_buffer_reg[23][1]  ( .D(\row2_buffer[24][1] ), .CK(clk), .Q(
        \row2_buffer[23][1] ) );
  DFFQXL \row2_buffer_reg[22][1]  ( .D(\row2_buffer[23][1] ), .CK(clk), .Q(
        \row2_buffer[22][1] ) );
  DFFQXL \row2_buffer_reg[21][1]  ( .D(\row2_buffer[22][1] ), .CK(clk), .Q(
        \row2_buffer[21][1] ) );
  DFFQXL \row2_buffer_reg[20][1]  ( .D(\row2_buffer[21][1] ), .CK(clk), .Q(
        \row2_buffer[20][1] ) );
  DFFQXL \row2_buffer_reg[19][1]  ( .D(\row2_buffer[20][1] ), .CK(clk), .Q(
        \row2_buffer[19][1] ) );
  DFFQXL \row2_buffer_reg[18][1]  ( .D(\row2_buffer[19][1] ), .CK(clk), .Q(
        \row2_buffer[18][1] ) );
  DFFQXL \row2_buffer_reg[17][1]  ( .D(\row2_buffer[18][1] ), .CK(clk), .Q(
        \row2_buffer[17][1] ) );
  DFFQXL \row2_buffer_reg[16][1]  ( .D(\row2_buffer[17][1] ), .CK(clk), .Q(
        \row2_buffer[16][1] ) );
  DFFQXL \row2_buffer_reg[15][1]  ( .D(\row2_buffer[16][1] ), .CK(clk), .Q(
        \row2_buffer[15][1] ) );
  DFFQXL \row2_buffer_reg[14][1]  ( .D(\row2_buffer[15][1] ), .CK(clk), .Q(
        \row2_buffer[14][1] ) );
  DFFQXL \row2_buffer_reg[13][1]  ( .D(\row2_buffer[14][1] ), .CK(clk), .Q(
        \row2_buffer[13][1] ) );
  DFFQXL \row2_buffer_reg[12][1]  ( .D(\row2_buffer[13][1] ), .CK(clk), .Q(
        \row2_buffer[12][1] ) );
  DFFQXL \row2_buffer_reg[11][1]  ( .D(\row2_buffer[12][1] ), .CK(clk), .Q(
        \row2_buffer[11][1] ) );
  DFFQXL \row2_buffer_reg[10][1]  ( .D(\row2_buffer[11][1] ), .CK(clk), .Q(
        \row2_buffer[10][1] ) );
  DFFQXL \row2_buffer_reg[9][1]  ( .D(\row2_buffer[10][1] ), .CK(clk), .Q(
        \row2_buffer[9][1] ) );
  DFFQXL \row2_buffer_reg[8][1]  ( .D(\row2_buffer[9][1] ), .CK(clk), .Q(
        \row2_buffer[8][1] ) );
  DFFQXL \row2_buffer_reg[7][1]  ( .D(\row2_buffer[8][1] ), .CK(clk), .Q(
        \row2_buffer[7][1] ) );
  DFFQXL \row2_buffer_reg[6][1]  ( .D(\row2_buffer[7][1] ), .CK(clk), .Q(
        \row2_buffer[6][1] ) );
  DFFQXL \row2_buffer_reg[5][1]  ( .D(\row2_buffer[6][1] ), .CK(clk), .Q(
        \row2_buffer[5][1] ) );
  DFFQXL \row2_buffer_reg[4][1]  ( .D(\row2_buffer[5][1] ), .CK(clk), .Q(
        \row2_buffer[4][1] ) );
  DFFQXL \row2_buffer_reg[3][1]  ( .D(\row2_buffer[4][1] ), .CK(clk), .Q(
        \row2_buffer[3][1] ) );
  DFFQXL \row1_buffer_reg[225][1]  ( .D(\row2_buffer[0][1] ), .CK(clk), .Q(
        \row1_buffer[225][1] ) );
  DFFQXL \row1_buffer_reg[224][1]  ( .D(\row1_buffer[225][1] ), .CK(clk), .Q(
        \row1_buffer[224][1] ) );
  DFFQXL \row1_buffer_reg[223][1]  ( .D(\row1_buffer[224][1] ), .CK(clk), .Q(
        \row1_buffer[223][1] ) );
  DFFQXL \row1_buffer_reg[222][1]  ( .D(\row1_buffer[223][1] ), .CK(clk), .Q(
        \row1_buffer[222][1] ) );
  DFFQXL \row1_buffer_reg[221][1]  ( .D(\row1_buffer[222][1] ), .CK(clk), .Q(
        \row1_buffer[221][1] ) );
  DFFQXL \row1_buffer_reg[220][1]  ( .D(\row1_buffer[221][1] ), .CK(clk), .Q(
        \row1_buffer[220][1] ) );
  DFFQXL \row1_buffer_reg[219][1]  ( .D(\row1_buffer[220][1] ), .CK(clk), .Q(
        \row1_buffer[219][1] ) );
  DFFQXL \row1_buffer_reg[218][1]  ( .D(\row1_buffer[219][1] ), .CK(clk), .Q(
        \row1_buffer[218][1] ) );
  DFFQXL \row1_buffer_reg[217][1]  ( .D(\row1_buffer[218][1] ), .CK(clk), .Q(
        \row1_buffer[217][1] ) );
  DFFQXL \row1_buffer_reg[216][1]  ( .D(\row1_buffer[217][1] ), .CK(clk), .Q(
        \row1_buffer[216][1] ) );
  DFFQXL \row1_buffer_reg[215][1]  ( .D(\row1_buffer[216][1] ), .CK(clk), .Q(
        \row1_buffer[215][1] ) );
  DFFQXL \row1_buffer_reg[214][1]  ( .D(\row1_buffer[215][1] ), .CK(clk), .Q(
        \row1_buffer[214][1] ) );
  DFFQXL \row1_buffer_reg[213][1]  ( .D(\row1_buffer[214][1] ), .CK(clk), .Q(
        \row1_buffer[213][1] ) );
  DFFQXL \row1_buffer_reg[212][1]  ( .D(\row1_buffer[213][1] ), .CK(clk), .Q(
        \row1_buffer[212][1] ) );
  DFFQXL \row1_buffer_reg[211][1]  ( .D(\row1_buffer[212][1] ), .CK(clk), .Q(
        \row1_buffer[211][1] ) );
  DFFQXL \row1_buffer_reg[210][1]  ( .D(\row1_buffer[211][1] ), .CK(clk), .Q(
        \row1_buffer[210][1] ) );
  DFFQXL \row1_buffer_reg[209][1]  ( .D(\row1_buffer[210][1] ), .CK(clk), .Q(
        \row1_buffer[209][1] ) );
  DFFQXL \row1_buffer_reg[208][1]  ( .D(\row1_buffer[209][1] ), .CK(clk), .Q(
        \row1_buffer[208][1] ) );
  DFFQXL \row1_buffer_reg[207][1]  ( .D(\row1_buffer[208][1] ), .CK(clk), .Q(
        \row1_buffer[207][1] ) );
  DFFQXL \row1_buffer_reg[206][1]  ( .D(\row1_buffer[207][1] ), .CK(clk), .Q(
        \row1_buffer[206][1] ) );
  DFFQXL \row1_buffer_reg[205][1]  ( .D(\row1_buffer[206][1] ), .CK(clk), .Q(
        \row1_buffer[205][1] ) );
  DFFQXL \row1_buffer_reg[204][1]  ( .D(\row1_buffer[205][1] ), .CK(clk), .Q(
        \row1_buffer[204][1] ) );
  DFFQXL \row1_buffer_reg[203][1]  ( .D(\row1_buffer[204][1] ), .CK(clk), .Q(
        \row1_buffer[203][1] ) );
  DFFQXL \row1_buffer_reg[202][1]  ( .D(\row1_buffer[203][1] ), .CK(clk), .Q(
        \row1_buffer[202][1] ) );
  DFFQXL \row1_buffer_reg[201][1]  ( .D(\row1_buffer[202][1] ), .CK(clk), .Q(
        \row1_buffer[201][1] ) );
  DFFQXL \row1_buffer_reg[200][1]  ( .D(\row1_buffer[201][1] ), .CK(clk), .Q(
        \row1_buffer[200][1] ) );
  DFFQXL \row1_buffer_reg[199][1]  ( .D(\row1_buffer[200][1] ), .CK(clk), .Q(
        \row1_buffer[199][1] ) );
  DFFQXL \row1_buffer_reg[198][1]  ( .D(\row1_buffer[199][1] ), .CK(clk), .Q(
        \row1_buffer[198][1] ) );
  DFFQXL \row1_buffer_reg[197][1]  ( .D(\row1_buffer[198][1] ), .CK(clk), .Q(
        \row1_buffer[197][1] ) );
  DFFQXL \row1_buffer_reg[196][1]  ( .D(\row1_buffer[197][1] ), .CK(clk), .Q(
        \row1_buffer[196][1] ) );
  DFFQXL \row1_buffer_reg[195][1]  ( .D(\row1_buffer[196][1] ), .CK(clk), .Q(
        \row1_buffer[195][1] ) );
  DFFQXL \row1_buffer_reg[194][1]  ( .D(\row1_buffer[195][1] ), .CK(clk), .Q(
        \row1_buffer[194][1] ) );
  DFFQXL \row1_buffer_reg[193][1]  ( .D(\row1_buffer[194][1] ), .CK(clk), .Q(
        \row1_buffer[193][1] ) );
  DFFQXL \row1_buffer_reg[192][1]  ( .D(\row1_buffer[193][1] ), .CK(clk), .Q(
        \row1_buffer[192][1] ) );
  DFFQXL \row1_buffer_reg[191][1]  ( .D(\row1_buffer[192][1] ), .CK(clk), .Q(
        \row1_buffer[191][1] ) );
  DFFQXL \row1_buffer_reg[190][1]  ( .D(\row1_buffer[191][1] ), .CK(clk), .Q(
        \row1_buffer[190][1] ) );
  DFFQXL \row1_buffer_reg[189][1]  ( .D(\row1_buffer[190][1] ), .CK(clk), .Q(
        \row1_buffer[189][1] ) );
  DFFQXL \row1_buffer_reg[188][1]  ( .D(\row1_buffer[189][1] ), .CK(clk), .Q(
        \row1_buffer[188][1] ) );
  DFFQXL \row1_buffer_reg[187][1]  ( .D(\row1_buffer[188][1] ), .CK(clk), .Q(
        \row1_buffer[187][1] ) );
  DFFQXL \row1_buffer_reg[186][1]  ( .D(\row1_buffer[187][1] ), .CK(clk), .Q(
        \row1_buffer[186][1] ) );
  DFFQXL \row1_buffer_reg[185][1]  ( .D(\row1_buffer[186][1] ), .CK(clk), .Q(
        \row1_buffer[185][1] ) );
  DFFQXL \row1_buffer_reg[184][1]  ( .D(\row1_buffer[185][1] ), .CK(clk), .Q(
        \row1_buffer[184][1] ) );
  DFFQXL \row1_buffer_reg[183][1]  ( .D(\row1_buffer[184][1] ), .CK(clk), .Q(
        \row1_buffer[183][1] ) );
  DFFQXL \row1_buffer_reg[182][1]  ( .D(\row1_buffer[183][1] ), .CK(clk), .Q(
        \row1_buffer[182][1] ) );
  DFFQXL \row1_buffer_reg[181][1]  ( .D(\row1_buffer[182][1] ), .CK(clk), .Q(
        \row1_buffer[181][1] ) );
  DFFQXL \row1_buffer_reg[180][1]  ( .D(\row1_buffer[181][1] ), .CK(clk), .Q(
        \row1_buffer[180][1] ) );
  DFFQXL \row1_buffer_reg[179][1]  ( .D(\row1_buffer[180][1] ), .CK(clk), .Q(
        \row1_buffer[179][1] ) );
  DFFQXL \row1_buffer_reg[178][1]  ( .D(\row1_buffer[179][1] ), .CK(clk), .Q(
        \row1_buffer[178][1] ) );
  DFFQXL \row1_buffer_reg[177][1]  ( .D(\row1_buffer[178][1] ), .CK(clk), .Q(
        \row1_buffer[177][1] ) );
  DFFQXL \row1_buffer_reg[176][1]  ( .D(\row1_buffer[177][1] ), .CK(clk), .Q(
        \row1_buffer[176][1] ) );
  DFFQXL \row1_buffer_reg[175][1]  ( .D(\row1_buffer[176][1] ), .CK(clk), .Q(
        \row1_buffer[175][1] ) );
  DFFQXL \row1_buffer_reg[174][1]  ( .D(\row1_buffer[175][1] ), .CK(clk), .Q(
        \row1_buffer[174][1] ) );
  DFFQXL \row1_buffer_reg[173][1]  ( .D(\row1_buffer[174][1] ), .CK(clk), .Q(
        \row1_buffer[173][1] ) );
  DFFQXL \row1_buffer_reg[172][1]  ( .D(\row1_buffer[173][1] ), .CK(clk), .Q(
        \row1_buffer[172][1] ) );
  DFFQXL \row1_buffer_reg[171][1]  ( .D(\row1_buffer[172][1] ), .CK(clk), .Q(
        \row1_buffer[171][1] ) );
  DFFQXL \row1_buffer_reg[170][1]  ( .D(\row1_buffer[171][1] ), .CK(clk), .Q(
        \row1_buffer[170][1] ) );
  DFFQXL \row1_buffer_reg[169][1]  ( .D(\row1_buffer[170][1] ), .CK(clk), .Q(
        \row1_buffer[169][1] ) );
  DFFQXL \row1_buffer_reg[168][1]  ( .D(\row1_buffer[169][1] ), .CK(clk), .Q(
        \row1_buffer[168][1] ) );
  DFFQXL \row1_buffer_reg[167][1]  ( .D(\row1_buffer[168][1] ), .CK(clk), .Q(
        \row1_buffer[167][1] ) );
  DFFQXL \row1_buffer_reg[166][1]  ( .D(\row1_buffer[167][1] ), .CK(clk), .Q(
        \row1_buffer[166][1] ) );
  DFFQXL \row1_buffer_reg[165][1]  ( .D(\row1_buffer[166][1] ), .CK(clk), .Q(
        \row1_buffer[165][1] ) );
  DFFQXL \row1_buffer_reg[164][1]  ( .D(\row1_buffer[165][1] ), .CK(clk), .Q(
        \row1_buffer[164][1] ) );
  DFFQXL \row1_buffer_reg[163][1]  ( .D(\row1_buffer[164][1] ), .CK(clk), .Q(
        \row1_buffer[163][1] ) );
  DFFQXL \row1_buffer_reg[162][1]  ( .D(\row1_buffer[163][1] ), .CK(clk), .Q(
        \row1_buffer[162][1] ) );
  DFFQXL \row1_buffer_reg[161][1]  ( .D(\row1_buffer[162][1] ), .CK(clk), .Q(
        \row1_buffer[161][1] ) );
  DFFQXL \row1_buffer_reg[160][1]  ( .D(\row1_buffer[161][1] ), .CK(clk), .Q(
        \row1_buffer[160][1] ) );
  DFFQXL \row1_buffer_reg[159][1]  ( .D(\row1_buffer[160][1] ), .CK(clk), .Q(
        \row1_buffer[159][1] ) );
  DFFQXL \row1_buffer_reg[158][1]  ( .D(\row1_buffer[159][1] ), .CK(clk), .Q(
        \row1_buffer[158][1] ) );
  DFFQXL \row1_buffer_reg[157][1]  ( .D(\row1_buffer[158][1] ), .CK(clk), .Q(
        \row1_buffer[157][1] ) );
  DFFQXL \row1_buffer_reg[156][1]  ( .D(\row1_buffer[157][1] ), .CK(clk), .Q(
        \row1_buffer[156][1] ) );
  DFFQXL \row1_buffer_reg[155][1]  ( .D(\row1_buffer[156][1] ), .CK(clk), .Q(
        \row1_buffer[155][1] ) );
  DFFQXL \row1_buffer_reg[154][1]  ( .D(\row1_buffer[155][1] ), .CK(clk), .Q(
        \row1_buffer[154][1] ) );
  DFFQXL \row1_buffer_reg[153][1]  ( .D(\row1_buffer[154][1] ), .CK(clk), .Q(
        \row1_buffer[153][1] ) );
  DFFQXL \row1_buffer_reg[152][1]  ( .D(\row1_buffer[153][1] ), .CK(clk), .Q(
        \row1_buffer[152][1] ) );
  DFFQXL \row1_buffer_reg[151][1]  ( .D(\row1_buffer[152][1] ), .CK(clk), .Q(
        \row1_buffer[151][1] ) );
  DFFQXL \row1_buffer_reg[150][1]  ( .D(\row1_buffer[151][1] ), .CK(clk), .Q(
        \row1_buffer[150][1] ) );
  DFFQXL \row1_buffer_reg[149][1]  ( .D(\row1_buffer[150][1] ), .CK(clk), .Q(
        \row1_buffer[149][1] ) );
  DFFQXL \row1_buffer_reg[148][1]  ( .D(\row1_buffer[149][1] ), .CK(clk), .Q(
        \row1_buffer[148][1] ) );
  DFFQXL \row1_buffer_reg[147][1]  ( .D(\row1_buffer[148][1] ), .CK(clk), .Q(
        \row1_buffer[147][1] ) );
  DFFQXL \row1_buffer_reg[146][1]  ( .D(\row1_buffer[147][1] ), .CK(clk), .Q(
        \row1_buffer[146][1] ) );
  DFFQXL \row1_buffer_reg[145][1]  ( .D(\row1_buffer[146][1] ), .CK(clk), .Q(
        \row1_buffer[145][1] ) );
  DFFQXL \row1_buffer_reg[144][1]  ( .D(\row1_buffer[145][1] ), .CK(clk), .Q(
        \row1_buffer[144][1] ) );
  DFFQXL \row1_buffer_reg[143][1]  ( .D(\row1_buffer[144][1] ), .CK(clk), .Q(
        \row1_buffer[143][1] ) );
  DFFQXL \row1_buffer_reg[142][1]  ( .D(\row1_buffer[143][1] ), .CK(clk), .Q(
        \row1_buffer[142][1] ) );
  DFFQXL \row1_buffer_reg[141][1]  ( .D(\row1_buffer[142][1] ), .CK(clk), .Q(
        \row1_buffer[141][1] ) );
  DFFQXL \row1_buffer_reg[140][1]  ( .D(\row1_buffer[141][1] ), .CK(clk), .Q(
        \row1_buffer[140][1] ) );
  DFFQXL \row1_buffer_reg[139][1]  ( .D(\row1_buffer[140][1] ), .CK(clk), .Q(
        \row1_buffer[139][1] ) );
  DFFQXL \row1_buffer_reg[138][1]  ( .D(\row1_buffer[139][1] ), .CK(clk), .Q(
        \row1_buffer[138][1] ) );
  DFFQXL \row1_buffer_reg[137][1]  ( .D(\row1_buffer[138][1] ), .CK(clk), .Q(
        \row1_buffer[137][1] ) );
  DFFQXL \row1_buffer_reg[136][1]  ( .D(\row1_buffer[137][1] ), .CK(clk), .Q(
        \row1_buffer[136][1] ) );
  DFFQXL \row1_buffer_reg[135][1]  ( .D(\row1_buffer[136][1] ), .CK(clk), .Q(
        \row1_buffer[135][1] ) );
  DFFQXL \row1_buffer_reg[134][1]  ( .D(\row1_buffer[135][1] ), .CK(clk), .Q(
        \row1_buffer[134][1] ) );
  DFFQXL \row1_buffer_reg[133][1]  ( .D(\row1_buffer[134][1] ), .CK(clk), .Q(
        \row1_buffer[133][1] ) );
  DFFQXL \row1_buffer_reg[132][1]  ( .D(\row1_buffer[133][1] ), .CK(clk), .Q(
        \row1_buffer[132][1] ) );
  DFFQXL \row1_buffer_reg[131][1]  ( .D(\row1_buffer[132][1] ), .CK(clk), .Q(
        \row1_buffer[131][1] ) );
  DFFQXL \row1_buffer_reg[130][1]  ( .D(\row1_buffer[131][1] ), .CK(clk), .Q(
        \row1_buffer[130][1] ) );
  DFFQXL \row1_buffer_reg[129][1]  ( .D(\row1_buffer[130][1] ), .CK(clk), .Q(
        \row1_buffer[129][1] ) );
  DFFQXL \row1_buffer_reg[128][1]  ( .D(\row1_buffer[129][1] ), .CK(clk), .Q(
        \row1_buffer[128][1] ) );
  DFFQXL \row1_buffer_reg[127][1]  ( .D(\row1_buffer[128][1] ), .CK(clk), .Q(
        \row1_buffer[127][1] ) );
  DFFQXL \row1_buffer_reg[126][1]  ( .D(\row1_buffer[127][1] ), .CK(clk), .Q(
        \row1_buffer[126][1] ) );
  DFFQXL \row1_buffer_reg[125][1]  ( .D(\row1_buffer[126][1] ), .CK(clk), .Q(
        \row1_buffer[125][1] ) );
  DFFQXL \row1_buffer_reg[124][1]  ( .D(\row1_buffer[125][1] ), .CK(clk), .Q(
        \row1_buffer[124][1] ) );
  DFFQXL \row1_buffer_reg[123][1]  ( .D(\row1_buffer[124][1] ), .CK(clk), .Q(
        \row1_buffer[123][1] ) );
  DFFQXL \row1_buffer_reg[122][1]  ( .D(\row1_buffer[123][1] ), .CK(clk), .Q(
        \row1_buffer[122][1] ) );
  DFFQXL \row1_buffer_reg[121][1]  ( .D(\row1_buffer[122][1] ), .CK(clk), .Q(
        \row1_buffer[121][1] ) );
  DFFQXL \row1_buffer_reg[120][1]  ( .D(\row1_buffer[121][1] ), .CK(clk), .Q(
        \row1_buffer[120][1] ) );
  DFFQXL \row1_buffer_reg[119][1]  ( .D(\row1_buffer[120][1] ), .CK(clk), .Q(
        \row1_buffer[119][1] ) );
  DFFQXL \row1_buffer_reg[118][1]  ( .D(\row1_buffer[119][1] ), .CK(clk), .Q(
        \row1_buffer[118][1] ) );
  DFFQXL \row1_buffer_reg[117][1]  ( .D(\row1_buffer[118][1] ), .CK(clk), .Q(
        \row1_buffer[117][1] ) );
  DFFQXL \row1_buffer_reg[116][1]  ( .D(\row1_buffer[117][1] ), .CK(clk), .Q(
        \row1_buffer[116][1] ) );
  DFFQXL \row1_buffer_reg[115][1]  ( .D(\row1_buffer[116][1] ), .CK(clk), .Q(
        \row1_buffer[115][1] ) );
  DFFQXL \row1_buffer_reg[114][1]  ( .D(\row1_buffer[115][1] ), .CK(clk), .Q(
        \row1_buffer[114][1] ) );
  DFFQXL \row1_buffer_reg[113][1]  ( .D(\row1_buffer[114][1] ), .CK(clk), .Q(
        \row1_buffer[113][1] ) );
  DFFQXL \row1_buffer_reg[112][1]  ( .D(\row1_buffer[113][1] ), .CK(clk), .Q(
        \row1_buffer[112][1] ) );
  DFFQXL \row1_buffer_reg[111][1]  ( .D(\row1_buffer[112][1] ), .CK(clk), .Q(
        \row1_buffer[111][1] ) );
  DFFQXL \row1_buffer_reg[110][1]  ( .D(\row1_buffer[111][1] ), .CK(clk), .Q(
        \row1_buffer[110][1] ) );
  DFFQXL \row1_buffer_reg[109][1]  ( .D(\row1_buffer[110][1] ), .CK(clk), .Q(
        \row1_buffer[109][1] ) );
  DFFQXL \row1_buffer_reg[108][1]  ( .D(\row1_buffer[109][1] ), .CK(clk), .Q(
        \row1_buffer[108][1] ) );
  DFFQXL \row1_buffer_reg[107][1]  ( .D(\row1_buffer[108][1] ), .CK(clk), .Q(
        \row1_buffer[107][1] ) );
  DFFQXL \row1_buffer_reg[106][1]  ( .D(\row1_buffer[107][1] ), .CK(clk), .Q(
        \row1_buffer[106][1] ) );
  DFFQXL \row1_buffer_reg[105][1]  ( .D(\row1_buffer[106][1] ), .CK(clk), .Q(
        \row1_buffer[105][1] ) );
  DFFQXL \row1_buffer_reg[104][1]  ( .D(\row1_buffer[105][1] ), .CK(clk), .Q(
        \row1_buffer[104][1] ) );
  DFFQXL \row1_buffer_reg[103][1]  ( .D(\row1_buffer[104][1] ), .CK(clk), .Q(
        \row1_buffer[103][1] ) );
  DFFQXL \row1_buffer_reg[102][1]  ( .D(\row1_buffer[103][1] ), .CK(clk), .Q(
        \row1_buffer[102][1] ) );
  DFFQXL \row1_buffer_reg[101][1]  ( .D(\row1_buffer[102][1] ), .CK(clk), .Q(
        \row1_buffer[101][1] ) );
  DFFQXL \row1_buffer_reg[100][1]  ( .D(\row1_buffer[101][1] ), .CK(clk), .Q(
        \row1_buffer[100][1] ) );
  DFFQXL \row1_buffer_reg[99][1]  ( .D(\row1_buffer[100][1] ), .CK(clk), .Q(
        \row1_buffer[99][1] ) );
  DFFQXL \row1_buffer_reg[98][1]  ( .D(\row1_buffer[99][1] ), .CK(clk), .Q(
        \row1_buffer[98][1] ) );
  DFFQXL \row1_buffer_reg[97][1]  ( .D(\row1_buffer[98][1] ), .CK(clk), .Q(
        \row1_buffer[97][1] ) );
  DFFQXL \row1_buffer_reg[96][1]  ( .D(\row1_buffer[97][1] ), .CK(clk), .Q(
        \row1_buffer[96][1] ) );
  DFFQXL \row1_buffer_reg[95][1]  ( .D(\row1_buffer[96][1] ), .CK(clk), .Q(
        \row1_buffer[95][1] ) );
  DFFQXL \row1_buffer_reg[94][1]  ( .D(\row1_buffer[95][1] ), .CK(clk), .Q(
        \row1_buffer[94][1] ) );
  DFFQXL \row1_buffer_reg[93][1]  ( .D(\row1_buffer[94][1] ), .CK(clk), .Q(
        \row1_buffer[93][1] ) );
  DFFQXL \row1_buffer_reg[92][1]  ( .D(\row1_buffer[93][1] ), .CK(clk), .Q(
        \row1_buffer[92][1] ) );
  DFFQXL \row1_buffer_reg[91][1]  ( .D(\row1_buffer[92][1] ), .CK(clk), .Q(
        \row1_buffer[91][1] ) );
  DFFQXL \row1_buffer_reg[90][1]  ( .D(\row1_buffer[91][1] ), .CK(clk), .Q(
        \row1_buffer[90][1] ) );
  DFFQXL \row1_buffer_reg[89][1]  ( .D(\row1_buffer[90][1] ), .CK(clk), .Q(
        \row1_buffer[89][1] ) );
  DFFQXL \row1_buffer_reg[88][1]  ( .D(\row1_buffer[89][1] ), .CK(clk), .Q(
        \row1_buffer[88][1] ) );
  DFFQXL \row1_buffer_reg[87][1]  ( .D(\row1_buffer[88][1] ), .CK(clk), .Q(
        \row1_buffer[87][1] ) );
  DFFQXL \row1_buffer_reg[86][1]  ( .D(\row1_buffer[87][1] ), .CK(clk), .Q(
        \row1_buffer[86][1] ) );
  DFFQXL \row1_buffer_reg[85][1]  ( .D(\row1_buffer[86][1] ), .CK(clk), .Q(
        \row1_buffer[85][1] ) );
  DFFQXL \row1_buffer_reg[84][1]  ( .D(\row1_buffer[85][1] ), .CK(clk), .Q(
        \row1_buffer[84][1] ) );
  DFFQXL \row1_buffer_reg[83][1]  ( .D(\row1_buffer[84][1] ), .CK(clk), .Q(
        \row1_buffer[83][1] ) );
  DFFQXL \row1_buffer_reg[82][1]  ( .D(\row1_buffer[83][1] ), .CK(clk), .Q(
        \row1_buffer[82][1] ) );
  DFFQXL \row1_buffer_reg[81][1]  ( .D(\row1_buffer[82][1] ), .CK(clk), .Q(
        \row1_buffer[81][1] ) );
  DFFQXL \row1_buffer_reg[80][1]  ( .D(\row1_buffer[81][1] ), .CK(clk), .Q(
        \row1_buffer[80][1] ) );
  DFFQXL \row1_buffer_reg[79][1]  ( .D(\row1_buffer[80][1] ), .CK(clk), .Q(
        \row1_buffer[79][1] ) );
  DFFQXL \row1_buffer_reg[78][1]  ( .D(\row1_buffer[79][1] ), .CK(clk), .Q(
        \row1_buffer[78][1] ) );
  DFFQXL \row1_buffer_reg[77][1]  ( .D(\row1_buffer[78][1] ), .CK(clk), .Q(
        \row1_buffer[77][1] ) );
  DFFQXL \row1_buffer_reg[76][1]  ( .D(\row1_buffer[77][1] ), .CK(clk), .Q(
        \row1_buffer[76][1] ) );
  DFFQXL \row1_buffer_reg[75][1]  ( .D(\row1_buffer[76][1] ), .CK(clk), .Q(
        \row1_buffer[75][1] ) );
  DFFQXL \row1_buffer_reg[74][1]  ( .D(\row1_buffer[75][1] ), .CK(clk), .Q(
        \row1_buffer[74][1] ) );
  DFFQXL \row1_buffer_reg[73][1]  ( .D(\row1_buffer[74][1] ), .CK(clk), .Q(
        \row1_buffer[73][1] ) );
  DFFQXL \row1_buffer_reg[72][1]  ( .D(\row1_buffer[73][1] ), .CK(clk), .Q(
        \row1_buffer[72][1] ) );
  DFFQXL \row1_buffer_reg[71][1]  ( .D(\row1_buffer[72][1] ), .CK(clk), .Q(
        \row1_buffer[71][1] ) );
  DFFQXL \row1_buffer_reg[70][1]  ( .D(\row1_buffer[71][1] ), .CK(clk), .Q(
        \row1_buffer[70][1] ) );
  DFFQXL \row1_buffer_reg[69][1]  ( .D(\row1_buffer[70][1] ), .CK(clk), .Q(
        \row1_buffer[69][1] ) );
  DFFQXL \row1_buffer_reg[68][1]  ( .D(\row1_buffer[69][1] ), .CK(clk), .Q(
        \row1_buffer[68][1] ) );
  DFFQXL \row1_buffer_reg[67][1]  ( .D(\row1_buffer[68][1] ), .CK(clk), .Q(
        \row1_buffer[67][1] ) );
  DFFQXL \row1_buffer_reg[66][1]  ( .D(\row1_buffer[67][1] ), .CK(clk), .Q(
        \row1_buffer[66][1] ) );
  DFFQXL \row1_buffer_reg[65][1]  ( .D(\row1_buffer[66][1] ), .CK(clk), .Q(
        \row1_buffer[65][1] ) );
  DFFQXL \row1_buffer_reg[64][1]  ( .D(\row1_buffer[65][1] ), .CK(clk), .Q(
        \row1_buffer[64][1] ) );
  DFFQXL \row1_buffer_reg[63][1]  ( .D(\row1_buffer[64][1] ), .CK(clk), .Q(
        \row1_buffer[63][1] ) );
  DFFQXL \row1_buffer_reg[62][1]  ( .D(\row1_buffer[63][1] ), .CK(clk), .Q(
        \row1_buffer[62][1] ) );
  DFFQXL \row1_buffer_reg[61][1]  ( .D(\row1_buffer[62][1] ), .CK(clk), .Q(
        \row1_buffer[61][1] ) );
  DFFQXL \row1_buffer_reg[60][1]  ( .D(\row1_buffer[61][1] ), .CK(clk), .Q(
        \row1_buffer[60][1] ) );
  DFFQXL \row1_buffer_reg[59][1]  ( .D(\row1_buffer[60][1] ), .CK(clk), .Q(
        \row1_buffer[59][1] ) );
  DFFQXL \row1_buffer_reg[58][1]  ( .D(\row1_buffer[59][1] ), .CK(clk), .Q(
        \row1_buffer[58][1] ) );
  DFFQXL \row1_buffer_reg[57][1]  ( .D(\row1_buffer[58][1] ), .CK(clk), .Q(
        \row1_buffer[57][1] ) );
  DFFQXL \row1_buffer_reg[56][1]  ( .D(\row1_buffer[57][1] ), .CK(clk), .Q(
        \row1_buffer[56][1] ) );
  DFFQXL \row1_buffer_reg[55][1]  ( .D(\row1_buffer[56][1] ), .CK(clk), .Q(
        \row1_buffer[55][1] ) );
  DFFQXL \row1_buffer_reg[54][1]  ( .D(\row1_buffer[55][1] ), .CK(clk), .Q(
        \row1_buffer[54][1] ) );
  DFFQXL \row1_buffer_reg[53][1]  ( .D(\row1_buffer[54][1] ), .CK(clk), .Q(
        \row1_buffer[53][1] ) );
  DFFQXL \row1_buffer_reg[52][1]  ( .D(\row1_buffer[53][1] ), .CK(clk), .Q(
        \row1_buffer[52][1] ) );
  DFFQXL \row1_buffer_reg[51][1]  ( .D(\row1_buffer[52][1] ), .CK(clk), .Q(
        \row1_buffer[51][1] ) );
  DFFQXL \row1_buffer_reg[50][1]  ( .D(\row1_buffer[51][1] ), .CK(clk), .Q(
        \row1_buffer[50][1] ) );
  DFFQXL \row1_buffer_reg[49][1]  ( .D(\row1_buffer[50][1] ), .CK(clk), .Q(
        \row1_buffer[49][1] ) );
  DFFQXL \row1_buffer_reg[48][1]  ( .D(\row1_buffer[49][1] ), .CK(clk), .Q(
        \row1_buffer[48][1] ) );
  DFFQXL \row1_buffer_reg[47][1]  ( .D(\row1_buffer[48][1] ), .CK(clk), .Q(
        \row1_buffer[47][1] ) );
  DFFQXL \row1_buffer_reg[46][1]  ( .D(\row1_buffer[47][1] ), .CK(clk), .Q(
        \row1_buffer[46][1] ) );
  DFFQXL \row1_buffer_reg[45][1]  ( .D(\row1_buffer[46][1] ), .CK(clk), .Q(
        \row1_buffer[45][1] ) );
  DFFQXL \row1_buffer_reg[44][1]  ( .D(\row1_buffer[45][1] ), .CK(clk), .Q(
        \row1_buffer[44][1] ) );
  DFFQXL \row1_buffer_reg[43][1]  ( .D(\row1_buffer[44][1] ), .CK(clk), .Q(
        \row1_buffer[43][1] ) );
  DFFQXL \row1_buffer_reg[42][1]  ( .D(\row1_buffer[43][1] ), .CK(clk), .Q(
        \row1_buffer[42][1] ) );
  DFFQXL \row1_buffer_reg[41][1]  ( .D(\row1_buffer[42][1] ), .CK(clk), .Q(
        \row1_buffer[41][1] ) );
  DFFQXL \row1_buffer_reg[40][1]  ( .D(\row1_buffer[41][1] ), .CK(clk), .Q(
        \row1_buffer[40][1] ) );
  DFFQXL \row1_buffer_reg[39][1]  ( .D(\row1_buffer[40][1] ), .CK(clk), .Q(
        \row1_buffer[39][1] ) );
  DFFQXL \row1_buffer_reg[38][1]  ( .D(\row1_buffer[39][1] ), .CK(clk), .Q(
        \row1_buffer[38][1] ) );
  DFFQXL \row1_buffer_reg[37][1]  ( .D(\row1_buffer[38][1] ), .CK(clk), .Q(
        \row1_buffer[37][1] ) );
  DFFQXL \row1_buffer_reg[36][1]  ( .D(\row1_buffer[37][1] ), .CK(clk), .Q(
        \row1_buffer[36][1] ) );
  DFFQXL \row1_buffer_reg[35][1]  ( .D(\row1_buffer[36][1] ), .CK(clk), .Q(
        \row1_buffer[35][1] ) );
  DFFQXL \row1_buffer_reg[34][1]  ( .D(\row1_buffer[35][1] ), .CK(clk), .Q(
        \row1_buffer[34][1] ) );
  DFFQXL \row1_buffer_reg[33][1]  ( .D(\row1_buffer[34][1] ), .CK(clk), .Q(
        \row1_buffer[33][1] ) );
  DFFQXL \row1_buffer_reg[32][1]  ( .D(\row1_buffer[33][1] ), .CK(clk), .Q(
        \row1_buffer[32][1] ) );
  DFFQXL \row1_buffer_reg[31][1]  ( .D(\row1_buffer[32][1] ), .CK(clk), .Q(
        \row1_buffer[31][1] ) );
  DFFQXL \row1_buffer_reg[30][1]  ( .D(\row1_buffer[31][1] ), .CK(clk), .Q(
        \row1_buffer[30][1] ) );
  DFFQXL \row1_buffer_reg[29][1]  ( .D(\row1_buffer[30][1] ), .CK(clk), .Q(
        \row1_buffer[29][1] ) );
  DFFQXL \row1_buffer_reg[28][1]  ( .D(\row1_buffer[29][1] ), .CK(clk), .Q(
        \row1_buffer[28][1] ) );
  DFFQXL \row1_buffer_reg[27][1]  ( .D(\row1_buffer[28][1] ), .CK(clk), .Q(
        \row1_buffer[27][1] ) );
  DFFQXL \row1_buffer_reg[26][1]  ( .D(\row1_buffer[27][1] ), .CK(clk), .Q(
        \row1_buffer[26][1] ) );
  DFFQXL \row1_buffer_reg[25][1]  ( .D(\row1_buffer[26][1] ), .CK(clk), .Q(
        \row1_buffer[25][1] ) );
  DFFQXL \row1_buffer_reg[24][1]  ( .D(\row1_buffer[25][1] ), .CK(clk), .Q(
        \row1_buffer[24][1] ) );
  DFFQXL \row1_buffer_reg[23][1]  ( .D(\row1_buffer[24][1] ), .CK(clk), .Q(
        \row1_buffer[23][1] ) );
  DFFQXL \row1_buffer_reg[22][1]  ( .D(\row1_buffer[23][1] ), .CK(clk), .Q(
        \row1_buffer[22][1] ) );
  DFFQXL \row1_buffer_reg[21][1]  ( .D(\row1_buffer[22][1] ), .CK(clk), .Q(
        \row1_buffer[21][1] ) );
  DFFQXL \row1_buffer_reg[20][1]  ( .D(\row1_buffer[21][1] ), .CK(clk), .Q(
        \row1_buffer[20][1] ) );
  DFFQXL \row1_buffer_reg[19][1]  ( .D(\row1_buffer[20][1] ), .CK(clk), .Q(
        \row1_buffer[19][1] ) );
  DFFQXL \row1_buffer_reg[18][1]  ( .D(\row1_buffer[19][1] ), .CK(clk), .Q(
        \row1_buffer[18][1] ) );
  DFFQXL \row1_buffer_reg[17][1]  ( .D(\row1_buffer[18][1] ), .CK(clk), .Q(
        \row1_buffer[17][1] ) );
  DFFQXL \row1_buffer_reg[16][1]  ( .D(\row1_buffer[17][1] ), .CK(clk), .Q(
        \row1_buffer[16][1] ) );
  DFFQXL \row1_buffer_reg[15][1]  ( .D(\row1_buffer[16][1] ), .CK(clk), .Q(
        \row1_buffer[15][1] ) );
  DFFQXL \row1_buffer_reg[14][1]  ( .D(\row1_buffer[15][1] ), .CK(clk), .Q(
        \row1_buffer[14][1] ) );
  DFFQXL \row1_buffer_reg[13][1]  ( .D(\row1_buffer[14][1] ), .CK(clk), .Q(
        \row1_buffer[13][1] ) );
  DFFQXL \row1_buffer_reg[12][1]  ( .D(\row1_buffer[13][1] ), .CK(clk), .Q(
        \row1_buffer[12][1] ) );
  DFFQXL \row1_buffer_reg[11][1]  ( .D(\row1_buffer[12][1] ), .CK(clk), .Q(
        \row1_buffer[11][1] ) );
  DFFQXL \row1_buffer_reg[10][1]  ( .D(\row1_buffer[11][1] ), .CK(clk), .Q(
        \row1_buffer[10][1] ) );
  DFFQXL \row1_buffer_reg[9][1]  ( .D(\row1_buffer[10][1] ), .CK(clk), .Q(
        \row1_buffer[9][1] ) );
  DFFQXL \row1_buffer_reg[8][1]  ( .D(\row1_buffer[9][1] ), .CK(clk), .Q(
        \row1_buffer[8][1] ) );
  DFFQXL \row1_buffer_reg[7][1]  ( .D(\row1_buffer[8][1] ), .CK(clk), .Q(
        \row1_buffer[7][1] ) );
  DFFQXL \row1_buffer_reg[6][1]  ( .D(\row1_buffer[7][1] ), .CK(clk), .Q(
        \row1_buffer[6][1] ) );
  DFFQXL \row1_buffer_reg[5][1]  ( .D(\row1_buffer[6][1] ), .CK(clk), .Q(
        \row1_buffer[5][1] ) );
  DFFQXL \row1_buffer_reg[4][1]  ( .D(\row1_buffer[5][1] ), .CK(clk), .Q(
        \row1_buffer[4][1] ) );
  DFFQXL \row1_buffer_reg[3][1]  ( .D(\row1_buffer[4][1] ), .CK(clk), .Q(
        \row1_buffer[3][1] ) );
  DFFQXL \row2_buffer_reg[225][0]  ( .D(\row3_buffer[0][0] ), .CK(clk), .Q(
        \row2_buffer[225][0] ) );
  DFFQXL \row2_buffer_reg[224][0]  ( .D(\row2_buffer[225][0] ), .CK(clk), .Q(
        \row2_buffer[224][0] ) );
  DFFQXL \row2_buffer_reg[223][0]  ( .D(\row2_buffer[224][0] ), .CK(clk), .Q(
        \row2_buffer[223][0] ) );
  DFFQXL \row2_buffer_reg[222][0]  ( .D(\row2_buffer[223][0] ), .CK(clk), .Q(
        \row2_buffer[222][0] ) );
  DFFQXL \row2_buffer_reg[221][0]  ( .D(\row2_buffer[222][0] ), .CK(clk), .Q(
        \row2_buffer[221][0] ) );
  DFFQXL \row2_buffer_reg[220][0]  ( .D(\row2_buffer[221][0] ), .CK(clk), .Q(
        \row2_buffer[220][0] ) );
  DFFQXL \row2_buffer_reg[219][0]  ( .D(\row2_buffer[220][0] ), .CK(clk), .Q(
        \row2_buffer[219][0] ) );
  DFFQXL \row2_buffer_reg[218][0]  ( .D(\row2_buffer[219][0] ), .CK(clk), .Q(
        \row2_buffer[218][0] ) );
  DFFQXL \row2_buffer_reg[217][0]  ( .D(\row2_buffer[218][0] ), .CK(clk), .Q(
        \row2_buffer[217][0] ) );
  DFFQXL \row2_buffer_reg[216][0]  ( .D(\row2_buffer[217][0] ), .CK(clk), .Q(
        \row2_buffer[216][0] ) );
  DFFQXL \row2_buffer_reg[215][0]  ( .D(\row2_buffer[216][0] ), .CK(clk), .Q(
        \row2_buffer[215][0] ) );
  DFFQXL \row2_buffer_reg[214][0]  ( .D(\row2_buffer[215][0] ), .CK(clk), .Q(
        \row2_buffer[214][0] ) );
  DFFQXL \row2_buffer_reg[213][0]  ( .D(\row2_buffer[214][0] ), .CK(clk), .Q(
        \row2_buffer[213][0] ) );
  DFFQXL \row2_buffer_reg[212][0]  ( .D(\row2_buffer[213][0] ), .CK(clk), .Q(
        \row2_buffer[212][0] ) );
  DFFQXL \row2_buffer_reg[211][0]  ( .D(\row2_buffer[212][0] ), .CK(clk), .Q(
        \row2_buffer[211][0] ) );
  DFFQXL \row2_buffer_reg[210][0]  ( .D(\row2_buffer[211][0] ), .CK(clk), .Q(
        \row2_buffer[210][0] ) );
  DFFQXL \row2_buffer_reg[209][0]  ( .D(\row2_buffer[210][0] ), .CK(clk), .Q(
        \row2_buffer[209][0] ) );
  DFFQXL \row2_buffer_reg[208][0]  ( .D(\row2_buffer[209][0] ), .CK(clk), .Q(
        \row2_buffer[208][0] ) );
  DFFQXL \row2_buffer_reg[207][0]  ( .D(\row2_buffer[208][0] ), .CK(clk), .Q(
        \row2_buffer[207][0] ) );
  DFFQXL \row2_buffer_reg[206][0]  ( .D(\row2_buffer[207][0] ), .CK(clk), .Q(
        \row2_buffer[206][0] ) );
  DFFQXL \row2_buffer_reg[205][0]  ( .D(\row2_buffer[206][0] ), .CK(clk), .Q(
        \row2_buffer[205][0] ) );
  DFFQXL \row2_buffer_reg[204][0]  ( .D(\row2_buffer[205][0] ), .CK(clk), .Q(
        \row2_buffer[204][0] ) );
  DFFQXL \row2_buffer_reg[203][0]  ( .D(\row2_buffer[204][0] ), .CK(clk), .Q(
        \row2_buffer[203][0] ) );
  DFFQXL \row2_buffer_reg[202][0]  ( .D(\row2_buffer[203][0] ), .CK(clk), .Q(
        \row2_buffer[202][0] ) );
  DFFQXL \row2_buffer_reg[201][0]  ( .D(\row2_buffer[202][0] ), .CK(clk), .Q(
        \row2_buffer[201][0] ) );
  DFFQXL \row2_buffer_reg[200][0]  ( .D(\row2_buffer[201][0] ), .CK(clk), .Q(
        \row2_buffer[200][0] ) );
  DFFQXL \row2_buffer_reg[199][0]  ( .D(\row2_buffer[200][0] ), .CK(clk), .Q(
        \row2_buffer[199][0] ) );
  DFFQXL \row2_buffer_reg[198][0]  ( .D(\row2_buffer[199][0] ), .CK(clk), .Q(
        \row2_buffer[198][0] ) );
  DFFQXL \row2_buffer_reg[197][0]  ( .D(\row2_buffer[198][0] ), .CK(clk), .Q(
        \row2_buffer[197][0] ) );
  DFFQXL \row2_buffer_reg[196][0]  ( .D(\row2_buffer[197][0] ), .CK(clk), .Q(
        \row2_buffer[196][0] ) );
  DFFQXL \row2_buffer_reg[195][0]  ( .D(\row2_buffer[196][0] ), .CK(clk), .Q(
        \row2_buffer[195][0] ) );
  DFFQXL \row2_buffer_reg[194][0]  ( .D(\row2_buffer[195][0] ), .CK(clk), .Q(
        \row2_buffer[194][0] ) );
  DFFQXL \row2_buffer_reg[193][0]  ( .D(\row2_buffer[194][0] ), .CK(clk), .Q(
        \row2_buffer[193][0] ) );
  DFFQXL \row2_buffer_reg[192][0]  ( .D(\row2_buffer[193][0] ), .CK(clk), .Q(
        \row2_buffer[192][0] ) );
  DFFQXL \row2_buffer_reg[191][0]  ( .D(\row2_buffer[192][0] ), .CK(clk), .Q(
        \row2_buffer[191][0] ) );
  DFFQXL \row2_buffer_reg[190][0]  ( .D(\row2_buffer[191][0] ), .CK(clk), .Q(
        \row2_buffer[190][0] ) );
  DFFQXL \row2_buffer_reg[189][0]  ( .D(\row2_buffer[190][0] ), .CK(clk), .Q(
        \row2_buffer[189][0] ) );
  DFFQXL \row2_buffer_reg[188][0]  ( .D(\row2_buffer[189][0] ), .CK(clk), .Q(
        \row2_buffer[188][0] ) );
  DFFQXL \row2_buffer_reg[187][0]  ( .D(\row2_buffer[188][0] ), .CK(clk), .Q(
        \row2_buffer[187][0] ) );
  DFFQXL \row2_buffer_reg[186][0]  ( .D(\row2_buffer[187][0] ), .CK(clk), .Q(
        \row2_buffer[186][0] ) );
  DFFQXL \row2_buffer_reg[185][0]  ( .D(\row2_buffer[186][0] ), .CK(clk), .Q(
        \row2_buffer[185][0] ) );
  DFFQXL \row2_buffer_reg[184][0]  ( .D(\row2_buffer[185][0] ), .CK(clk), .Q(
        \row2_buffer[184][0] ) );
  DFFQXL \row2_buffer_reg[183][0]  ( .D(\row2_buffer[184][0] ), .CK(clk), .Q(
        \row2_buffer[183][0] ) );
  DFFQXL \row2_buffer_reg[182][0]  ( .D(\row2_buffer[183][0] ), .CK(clk), .Q(
        \row2_buffer[182][0] ) );
  DFFQXL \row2_buffer_reg[181][0]  ( .D(\row2_buffer[182][0] ), .CK(clk), .Q(
        \row2_buffer[181][0] ) );
  DFFQXL \row2_buffer_reg[180][0]  ( .D(\row2_buffer[181][0] ), .CK(clk), .Q(
        \row2_buffer[180][0] ) );
  DFFQXL \row2_buffer_reg[179][0]  ( .D(\row2_buffer[180][0] ), .CK(clk), .Q(
        \row2_buffer[179][0] ) );
  DFFQXL \row2_buffer_reg[178][0]  ( .D(\row2_buffer[179][0] ), .CK(clk), .Q(
        \row2_buffer[178][0] ) );
  DFFQXL \row2_buffer_reg[177][0]  ( .D(\row2_buffer[178][0] ), .CK(clk), .Q(
        \row2_buffer[177][0] ) );
  DFFQXL \row2_buffer_reg[176][0]  ( .D(\row2_buffer[177][0] ), .CK(clk), .Q(
        \row2_buffer[176][0] ) );
  DFFQXL \row2_buffer_reg[175][0]  ( .D(\row2_buffer[176][0] ), .CK(clk), .Q(
        \row2_buffer[175][0] ) );
  DFFQXL \row2_buffer_reg[174][0]  ( .D(\row2_buffer[175][0] ), .CK(clk), .Q(
        \row2_buffer[174][0] ) );
  DFFQXL \row2_buffer_reg[173][0]  ( .D(\row2_buffer[174][0] ), .CK(clk), .Q(
        \row2_buffer[173][0] ) );
  DFFQXL \row2_buffer_reg[172][0]  ( .D(\row2_buffer[173][0] ), .CK(clk), .Q(
        \row2_buffer[172][0] ) );
  DFFQXL \row2_buffer_reg[171][0]  ( .D(\row2_buffer[172][0] ), .CK(clk), .Q(
        \row2_buffer[171][0] ) );
  DFFQXL \row2_buffer_reg[170][0]  ( .D(\row2_buffer[171][0] ), .CK(clk), .Q(
        \row2_buffer[170][0] ) );
  DFFQXL \row2_buffer_reg[169][0]  ( .D(\row2_buffer[170][0] ), .CK(clk), .Q(
        \row2_buffer[169][0] ) );
  DFFQXL \row2_buffer_reg[168][0]  ( .D(\row2_buffer[169][0] ), .CK(clk), .Q(
        \row2_buffer[168][0] ) );
  DFFQXL \row2_buffer_reg[167][0]  ( .D(\row2_buffer[168][0] ), .CK(clk), .Q(
        \row2_buffer[167][0] ) );
  DFFQXL \row2_buffer_reg[166][0]  ( .D(\row2_buffer[167][0] ), .CK(clk), .Q(
        \row2_buffer[166][0] ) );
  DFFQXL \row2_buffer_reg[165][0]  ( .D(\row2_buffer[166][0] ), .CK(clk), .Q(
        \row2_buffer[165][0] ) );
  DFFQXL \row2_buffer_reg[164][0]  ( .D(\row2_buffer[165][0] ), .CK(clk), .Q(
        \row2_buffer[164][0] ) );
  DFFQXL \row2_buffer_reg[163][0]  ( .D(\row2_buffer[164][0] ), .CK(clk), .Q(
        \row2_buffer[163][0] ) );
  DFFQXL \row2_buffer_reg[162][0]  ( .D(\row2_buffer[163][0] ), .CK(clk), .Q(
        \row2_buffer[162][0] ) );
  DFFQXL \row2_buffer_reg[161][0]  ( .D(\row2_buffer[162][0] ), .CK(clk), .Q(
        \row2_buffer[161][0] ) );
  DFFQXL \row2_buffer_reg[160][0]  ( .D(\row2_buffer[161][0] ), .CK(clk), .Q(
        \row2_buffer[160][0] ) );
  DFFQXL \row2_buffer_reg[159][0]  ( .D(\row2_buffer[160][0] ), .CK(clk), .Q(
        \row2_buffer[159][0] ) );
  DFFQXL \row2_buffer_reg[158][0]  ( .D(\row2_buffer[159][0] ), .CK(clk), .Q(
        \row2_buffer[158][0] ) );
  DFFQXL \row2_buffer_reg[157][0]  ( .D(\row2_buffer[158][0] ), .CK(clk), .Q(
        \row2_buffer[157][0] ) );
  DFFQXL \row2_buffer_reg[156][0]  ( .D(\row2_buffer[157][0] ), .CK(clk), .Q(
        \row2_buffer[156][0] ) );
  DFFQXL \row2_buffer_reg[155][0]  ( .D(\row2_buffer[156][0] ), .CK(clk), .Q(
        \row2_buffer[155][0] ) );
  DFFQXL \row2_buffer_reg[154][0]  ( .D(\row2_buffer[155][0] ), .CK(clk), .Q(
        \row2_buffer[154][0] ) );
  DFFQXL \row2_buffer_reg[153][0]  ( .D(\row2_buffer[154][0] ), .CK(clk), .Q(
        \row2_buffer[153][0] ) );
  DFFQXL \row2_buffer_reg[152][0]  ( .D(\row2_buffer[153][0] ), .CK(clk), .Q(
        \row2_buffer[152][0] ) );
  DFFQXL \row2_buffer_reg[151][0]  ( .D(\row2_buffer[152][0] ), .CK(clk), .Q(
        \row2_buffer[151][0] ) );
  DFFQXL \row2_buffer_reg[150][0]  ( .D(\row2_buffer[151][0] ), .CK(clk), .Q(
        \row2_buffer[150][0] ) );
  DFFQXL \row2_buffer_reg[149][0]  ( .D(\row2_buffer[150][0] ), .CK(clk), .Q(
        \row2_buffer[149][0] ) );
  DFFQXL \row2_buffer_reg[148][0]  ( .D(\row2_buffer[149][0] ), .CK(clk), .Q(
        \row2_buffer[148][0] ) );
  DFFQXL \row2_buffer_reg[147][0]  ( .D(\row2_buffer[148][0] ), .CK(clk), .Q(
        \row2_buffer[147][0] ) );
  DFFQXL \row2_buffer_reg[146][0]  ( .D(\row2_buffer[147][0] ), .CK(clk), .Q(
        \row2_buffer[146][0] ) );
  DFFQXL \row2_buffer_reg[145][0]  ( .D(\row2_buffer[146][0] ), .CK(clk), .Q(
        \row2_buffer[145][0] ) );
  DFFQXL \row2_buffer_reg[144][0]  ( .D(\row2_buffer[145][0] ), .CK(clk), .Q(
        \row2_buffer[144][0] ) );
  DFFQXL \row2_buffer_reg[143][0]  ( .D(\row2_buffer[144][0] ), .CK(clk), .Q(
        \row2_buffer[143][0] ) );
  DFFQXL \row2_buffer_reg[142][0]  ( .D(\row2_buffer[143][0] ), .CK(clk), .Q(
        \row2_buffer[142][0] ) );
  DFFQXL \row2_buffer_reg[141][0]  ( .D(\row2_buffer[142][0] ), .CK(clk), .Q(
        \row2_buffer[141][0] ) );
  DFFQXL \row2_buffer_reg[140][0]  ( .D(\row2_buffer[141][0] ), .CK(clk), .Q(
        \row2_buffer[140][0] ) );
  DFFQXL \row2_buffer_reg[139][0]  ( .D(\row2_buffer[140][0] ), .CK(clk), .Q(
        \row2_buffer[139][0] ) );
  DFFQXL \row2_buffer_reg[138][0]  ( .D(\row2_buffer[139][0] ), .CK(clk), .Q(
        \row2_buffer[138][0] ) );
  DFFQXL \row2_buffer_reg[137][0]  ( .D(\row2_buffer[138][0] ), .CK(clk), .Q(
        \row2_buffer[137][0] ) );
  DFFQXL \row2_buffer_reg[136][0]  ( .D(\row2_buffer[137][0] ), .CK(clk), .Q(
        \row2_buffer[136][0] ) );
  DFFQXL \row2_buffer_reg[135][0]  ( .D(\row2_buffer[136][0] ), .CK(clk), .Q(
        \row2_buffer[135][0] ) );
  DFFQXL \row2_buffer_reg[134][0]  ( .D(\row2_buffer[135][0] ), .CK(clk), .Q(
        \row2_buffer[134][0] ) );
  DFFQXL \row2_buffer_reg[133][0]  ( .D(\row2_buffer[134][0] ), .CK(clk), .Q(
        \row2_buffer[133][0] ) );
  DFFQXL \row2_buffer_reg[132][0]  ( .D(\row2_buffer[133][0] ), .CK(clk), .Q(
        \row2_buffer[132][0] ) );
  DFFQXL \row2_buffer_reg[131][0]  ( .D(\row2_buffer[132][0] ), .CK(clk), .Q(
        \row2_buffer[131][0] ) );
  DFFQXL \row2_buffer_reg[130][0]  ( .D(\row2_buffer[131][0] ), .CK(clk), .Q(
        \row2_buffer[130][0] ) );
  DFFQXL \row2_buffer_reg[129][0]  ( .D(\row2_buffer[130][0] ), .CK(clk), .Q(
        \row2_buffer[129][0] ) );
  DFFQXL \row2_buffer_reg[128][0]  ( .D(\row2_buffer[129][0] ), .CK(clk), .Q(
        \row2_buffer[128][0] ) );
  DFFQXL \row2_buffer_reg[127][0]  ( .D(\row2_buffer[128][0] ), .CK(clk), .Q(
        \row2_buffer[127][0] ) );
  DFFQXL \row2_buffer_reg[126][0]  ( .D(\row2_buffer[127][0] ), .CK(clk), .Q(
        \row2_buffer[126][0] ) );
  DFFQXL \row2_buffer_reg[125][0]  ( .D(\row2_buffer[126][0] ), .CK(clk), .Q(
        \row2_buffer[125][0] ) );
  DFFQXL \row2_buffer_reg[124][0]  ( .D(\row2_buffer[125][0] ), .CK(clk), .Q(
        \row2_buffer[124][0] ) );
  DFFQXL \row2_buffer_reg[123][0]  ( .D(\row2_buffer[124][0] ), .CK(clk), .Q(
        \row2_buffer[123][0] ) );
  DFFQXL \row2_buffer_reg[122][0]  ( .D(\row2_buffer[123][0] ), .CK(clk), .Q(
        \row2_buffer[122][0] ) );
  DFFQXL \row2_buffer_reg[121][0]  ( .D(\row2_buffer[122][0] ), .CK(clk), .Q(
        \row2_buffer[121][0] ) );
  DFFQXL \row2_buffer_reg[120][0]  ( .D(\row2_buffer[121][0] ), .CK(clk), .Q(
        \row2_buffer[120][0] ) );
  DFFQXL \row2_buffer_reg[119][0]  ( .D(\row2_buffer[120][0] ), .CK(clk), .Q(
        \row2_buffer[119][0] ) );
  DFFQXL \row2_buffer_reg[118][0]  ( .D(\row2_buffer[119][0] ), .CK(clk), .Q(
        \row2_buffer[118][0] ) );
  DFFQXL \row2_buffer_reg[117][0]  ( .D(\row2_buffer[118][0] ), .CK(clk), .Q(
        \row2_buffer[117][0] ) );
  DFFQXL \row2_buffer_reg[116][0]  ( .D(\row2_buffer[117][0] ), .CK(clk), .Q(
        \row2_buffer[116][0] ) );
  DFFQXL \row2_buffer_reg[115][0]  ( .D(\row2_buffer[116][0] ), .CK(clk), .Q(
        \row2_buffer[115][0] ) );
  DFFQXL \row2_buffer_reg[114][0]  ( .D(\row2_buffer[115][0] ), .CK(clk), .Q(
        \row2_buffer[114][0] ) );
  DFFQXL \row2_buffer_reg[113][0]  ( .D(\row2_buffer[114][0] ), .CK(clk), .Q(
        \row2_buffer[113][0] ) );
  DFFQXL \row2_buffer_reg[112][0]  ( .D(\row2_buffer[113][0] ), .CK(clk), .Q(
        \row2_buffer[112][0] ) );
  DFFQXL \row2_buffer_reg[111][0]  ( .D(\row2_buffer[112][0] ), .CK(clk), .Q(
        \row2_buffer[111][0] ) );
  DFFQXL \row2_buffer_reg[110][0]  ( .D(\row2_buffer[111][0] ), .CK(clk), .Q(
        \row2_buffer[110][0] ) );
  DFFQXL \row2_buffer_reg[109][0]  ( .D(\row2_buffer[110][0] ), .CK(clk), .Q(
        \row2_buffer[109][0] ) );
  DFFQXL \row2_buffer_reg[108][0]  ( .D(\row2_buffer[109][0] ), .CK(clk), .Q(
        \row2_buffer[108][0] ) );
  DFFQXL \row2_buffer_reg[107][0]  ( .D(\row2_buffer[108][0] ), .CK(clk), .Q(
        \row2_buffer[107][0] ) );
  DFFQXL \row2_buffer_reg[106][0]  ( .D(\row2_buffer[107][0] ), .CK(clk), .Q(
        \row2_buffer[106][0] ) );
  DFFQXL \row2_buffer_reg[105][0]  ( .D(\row2_buffer[106][0] ), .CK(clk), .Q(
        \row2_buffer[105][0] ) );
  DFFQXL \row2_buffer_reg[104][0]  ( .D(\row2_buffer[105][0] ), .CK(clk), .Q(
        \row2_buffer[104][0] ) );
  DFFQXL \row2_buffer_reg[103][0]  ( .D(\row2_buffer[104][0] ), .CK(clk), .Q(
        \row2_buffer[103][0] ) );
  DFFQXL \row2_buffer_reg[102][0]  ( .D(\row2_buffer[103][0] ), .CK(clk), .Q(
        \row2_buffer[102][0] ) );
  DFFQXL \row2_buffer_reg[101][0]  ( .D(\row2_buffer[102][0] ), .CK(clk), .Q(
        \row2_buffer[101][0] ) );
  DFFQXL \row2_buffer_reg[100][0]  ( .D(\row2_buffer[101][0] ), .CK(clk), .Q(
        \row2_buffer[100][0] ) );
  DFFQXL \row2_buffer_reg[99][0]  ( .D(\row2_buffer[100][0] ), .CK(clk), .Q(
        \row2_buffer[99][0] ) );
  DFFQXL \row2_buffer_reg[98][0]  ( .D(\row2_buffer[99][0] ), .CK(clk), .Q(
        \row2_buffer[98][0] ) );
  DFFQXL \row2_buffer_reg[97][0]  ( .D(\row2_buffer[98][0] ), .CK(clk), .Q(
        \row2_buffer[97][0] ) );
  DFFQXL \row2_buffer_reg[96][0]  ( .D(\row2_buffer[97][0] ), .CK(clk), .Q(
        \row2_buffer[96][0] ) );
  DFFQXL \row2_buffer_reg[95][0]  ( .D(\row2_buffer[96][0] ), .CK(clk), .Q(
        \row2_buffer[95][0] ) );
  DFFQXL \row2_buffer_reg[94][0]  ( .D(\row2_buffer[95][0] ), .CK(clk), .Q(
        \row2_buffer[94][0] ) );
  DFFQXL \row2_buffer_reg[93][0]  ( .D(\row2_buffer[94][0] ), .CK(clk), .Q(
        \row2_buffer[93][0] ) );
  DFFQXL \row2_buffer_reg[92][0]  ( .D(\row2_buffer[93][0] ), .CK(clk), .Q(
        \row2_buffer[92][0] ) );
  DFFQXL \row2_buffer_reg[91][0]  ( .D(\row2_buffer[92][0] ), .CK(clk), .Q(
        \row2_buffer[91][0] ) );
  DFFQXL \row2_buffer_reg[90][0]  ( .D(\row2_buffer[91][0] ), .CK(clk), .Q(
        \row2_buffer[90][0] ) );
  DFFQXL \row2_buffer_reg[89][0]  ( .D(\row2_buffer[90][0] ), .CK(clk), .Q(
        \row2_buffer[89][0] ) );
  DFFQXL \row2_buffer_reg[88][0]  ( .D(\row2_buffer[89][0] ), .CK(clk), .Q(
        \row2_buffer[88][0] ) );
  DFFQXL \row2_buffer_reg[87][0]  ( .D(\row2_buffer[88][0] ), .CK(clk), .Q(
        \row2_buffer[87][0] ) );
  DFFQXL \row2_buffer_reg[86][0]  ( .D(\row2_buffer[87][0] ), .CK(clk), .Q(
        \row2_buffer[86][0] ) );
  DFFQXL \row2_buffer_reg[85][0]  ( .D(\row2_buffer[86][0] ), .CK(clk), .Q(
        \row2_buffer[85][0] ) );
  DFFQXL \row2_buffer_reg[84][0]  ( .D(\row2_buffer[85][0] ), .CK(clk), .Q(
        \row2_buffer[84][0] ) );
  DFFQXL \row2_buffer_reg[83][0]  ( .D(\row2_buffer[84][0] ), .CK(clk), .Q(
        \row2_buffer[83][0] ) );
  DFFQXL \row2_buffer_reg[82][0]  ( .D(\row2_buffer[83][0] ), .CK(clk), .Q(
        \row2_buffer[82][0] ) );
  DFFQXL \row2_buffer_reg[81][0]  ( .D(\row2_buffer[82][0] ), .CK(clk), .Q(
        \row2_buffer[81][0] ) );
  DFFQXL \row2_buffer_reg[80][0]  ( .D(\row2_buffer[81][0] ), .CK(clk), .Q(
        \row2_buffer[80][0] ) );
  DFFQXL \row2_buffer_reg[79][0]  ( .D(\row2_buffer[80][0] ), .CK(clk), .Q(
        \row2_buffer[79][0] ) );
  DFFQXL \row2_buffer_reg[78][0]  ( .D(\row2_buffer[79][0] ), .CK(clk), .Q(
        \row2_buffer[78][0] ) );
  DFFQXL \row2_buffer_reg[77][0]  ( .D(\row2_buffer[78][0] ), .CK(clk), .Q(
        \row2_buffer[77][0] ) );
  DFFQXL \row2_buffer_reg[76][0]  ( .D(\row2_buffer[77][0] ), .CK(clk), .Q(
        \row2_buffer[76][0] ) );
  DFFQXL \row2_buffer_reg[75][0]  ( .D(\row2_buffer[76][0] ), .CK(clk), .Q(
        \row2_buffer[75][0] ) );
  DFFQXL \row2_buffer_reg[74][0]  ( .D(\row2_buffer[75][0] ), .CK(clk), .Q(
        \row2_buffer[74][0] ) );
  DFFQXL \row2_buffer_reg[73][0]  ( .D(\row2_buffer[74][0] ), .CK(clk), .Q(
        \row2_buffer[73][0] ) );
  DFFQXL \row2_buffer_reg[72][0]  ( .D(\row2_buffer[73][0] ), .CK(clk), .Q(
        \row2_buffer[72][0] ) );
  DFFQXL \row2_buffer_reg[71][0]  ( .D(\row2_buffer[72][0] ), .CK(clk), .Q(
        \row2_buffer[71][0] ) );
  DFFQXL \row2_buffer_reg[70][0]  ( .D(\row2_buffer[71][0] ), .CK(clk), .Q(
        \row2_buffer[70][0] ) );
  DFFQXL \row2_buffer_reg[69][0]  ( .D(\row2_buffer[70][0] ), .CK(clk), .Q(
        \row2_buffer[69][0] ) );
  DFFQXL \row2_buffer_reg[68][0]  ( .D(\row2_buffer[69][0] ), .CK(clk), .Q(
        \row2_buffer[68][0] ) );
  DFFQXL \row2_buffer_reg[67][0]  ( .D(\row2_buffer[68][0] ), .CK(clk), .Q(
        \row2_buffer[67][0] ) );
  DFFQXL \row2_buffer_reg[66][0]  ( .D(\row2_buffer[67][0] ), .CK(clk), .Q(
        \row2_buffer[66][0] ) );
  DFFQXL \row2_buffer_reg[65][0]  ( .D(\row2_buffer[66][0] ), .CK(clk), .Q(
        \row2_buffer[65][0] ) );
  DFFQXL \row2_buffer_reg[64][0]  ( .D(\row2_buffer[65][0] ), .CK(clk), .Q(
        \row2_buffer[64][0] ) );
  DFFQXL \row2_buffer_reg[63][0]  ( .D(\row2_buffer[64][0] ), .CK(clk), .Q(
        \row2_buffer[63][0] ) );
  DFFQXL \row2_buffer_reg[62][0]  ( .D(\row2_buffer[63][0] ), .CK(clk), .Q(
        \row2_buffer[62][0] ) );
  DFFQXL \row2_buffer_reg[61][0]  ( .D(\row2_buffer[62][0] ), .CK(clk), .Q(
        \row2_buffer[61][0] ) );
  DFFQXL \row2_buffer_reg[60][0]  ( .D(\row2_buffer[61][0] ), .CK(clk), .Q(
        \row2_buffer[60][0] ) );
  DFFQXL \row2_buffer_reg[59][0]  ( .D(\row2_buffer[60][0] ), .CK(clk), .Q(
        \row2_buffer[59][0] ) );
  DFFQXL \row2_buffer_reg[58][0]  ( .D(\row2_buffer[59][0] ), .CK(clk), .Q(
        \row2_buffer[58][0] ) );
  DFFQXL \row2_buffer_reg[57][0]  ( .D(\row2_buffer[58][0] ), .CK(clk), .Q(
        \row2_buffer[57][0] ) );
  DFFQXL \row2_buffer_reg[56][0]  ( .D(\row2_buffer[57][0] ), .CK(clk), .Q(
        \row2_buffer[56][0] ) );
  DFFQXL \row2_buffer_reg[55][0]  ( .D(\row2_buffer[56][0] ), .CK(clk), .Q(
        \row2_buffer[55][0] ) );
  DFFQXL \row2_buffer_reg[54][0]  ( .D(\row2_buffer[55][0] ), .CK(clk), .Q(
        \row2_buffer[54][0] ) );
  DFFQXL \row2_buffer_reg[53][0]  ( .D(\row2_buffer[54][0] ), .CK(clk), .Q(
        \row2_buffer[53][0] ) );
  DFFQXL \row2_buffer_reg[52][0]  ( .D(\row2_buffer[53][0] ), .CK(clk), .Q(
        \row2_buffer[52][0] ) );
  DFFQXL \row2_buffer_reg[51][0]  ( .D(\row2_buffer[52][0] ), .CK(clk), .Q(
        \row2_buffer[51][0] ) );
  DFFQXL \row2_buffer_reg[50][0]  ( .D(\row2_buffer[51][0] ), .CK(clk), .Q(
        \row2_buffer[50][0] ) );
  DFFQXL \row2_buffer_reg[49][0]  ( .D(\row2_buffer[50][0] ), .CK(clk), .Q(
        \row2_buffer[49][0] ) );
  DFFQXL \row2_buffer_reg[48][0]  ( .D(\row2_buffer[49][0] ), .CK(clk), .Q(
        \row2_buffer[48][0] ) );
  DFFQXL \row2_buffer_reg[47][0]  ( .D(\row2_buffer[48][0] ), .CK(clk), .Q(
        \row2_buffer[47][0] ) );
  DFFQXL \row2_buffer_reg[46][0]  ( .D(\row2_buffer[47][0] ), .CK(clk), .Q(
        \row2_buffer[46][0] ) );
  DFFQXL \row2_buffer_reg[45][0]  ( .D(\row2_buffer[46][0] ), .CK(clk), .Q(
        \row2_buffer[45][0] ) );
  DFFQXL \row2_buffer_reg[44][0]  ( .D(\row2_buffer[45][0] ), .CK(clk), .Q(
        \row2_buffer[44][0] ) );
  DFFQXL \row2_buffer_reg[43][0]  ( .D(\row2_buffer[44][0] ), .CK(clk), .Q(
        \row2_buffer[43][0] ) );
  DFFQXL \row2_buffer_reg[42][0]  ( .D(\row2_buffer[43][0] ), .CK(clk), .Q(
        \row2_buffer[42][0] ) );
  DFFQXL \row2_buffer_reg[41][0]  ( .D(\row2_buffer[42][0] ), .CK(clk), .Q(
        \row2_buffer[41][0] ) );
  DFFQXL \row2_buffer_reg[40][0]  ( .D(\row2_buffer[41][0] ), .CK(clk), .Q(
        \row2_buffer[40][0] ) );
  DFFQXL \row2_buffer_reg[39][0]  ( .D(\row2_buffer[40][0] ), .CK(clk), .Q(
        \row2_buffer[39][0] ) );
  DFFQXL \row2_buffer_reg[38][0]  ( .D(\row2_buffer[39][0] ), .CK(clk), .Q(
        \row2_buffer[38][0] ) );
  DFFQXL \row2_buffer_reg[37][0]  ( .D(\row2_buffer[38][0] ), .CK(clk), .Q(
        \row2_buffer[37][0] ) );
  DFFQXL \row2_buffer_reg[36][0]  ( .D(\row2_buffer[37][0] ), .CK(clk), .Q(
        \row2_buffer[36][0] ) );
  DFFQXL \row2_buffer_reg[35][0]  ( .D(\row2_buffer[36][0] ), .CK(clk), .Q(
        \row2_buffer[35][0] ) );
  DFFQXL \row2_buffer_reg[34][0]  ( .D(\row2_buffer[35][0] ), .CK(clk), .Q(
        \row2_buffer[34][0] ) );
  DFFQXL \row2_buffer_reg[33][0]  ( .D(\row2_buffer[34][0] ), .CK(clk), .Q(
        \row2_buffer[33][0] ) );
  DFFQXL \row2_buffer_reg[32][0]  ( .D(\row2_buffer[33][0] ), .CK(clk), .Q(
        \row2_buffer[32][0] ) );
  DFFQXL \row2_buffer_reg[31][0]  ( .D(\row2_buffer[32][0] ), .CK(clk), .Q(
        \row2_buffer[31][0] ) );
  DFFQXL \row2_buffer_reg[30][0]  ( .D(\row2_buffer[31][0] ), .CK(clk), .Q(
        \row2_buffer[30][0] ) );
  DFFQXL \row2_buffer_reg[29][0]  ( .D(\row2_buffer[30][0] ), .CK(clk), .Q(
        \row2_buffer[29][0] ) );
  DFFQXL \row2_buffer_reg[28][0]  ( .D(\row2_buffer[29][0] ), .CK(clk), .Q(
        \row2_buffer[28][0] ) );
  DFFQXL \row2_buffer_reg[27][0]  ( .D(\row2_buffer[28][0] ), .CK(clk), .Q(
        \row2_buffer[27][0] ) );
  DFFQXL \row2_buffer_reg[26][0]  ( .D(\row2_buffer[27][0] ), .CK(clk), .Q(
        \row2_buffer[26][0] ) );
  DFFQXL \row2_buffer_reg[25][0]  ( .D(\row2_buffer[26][0] ), .CK(clk), .Q(
        \row2_buffer[25][0] ) );
  DFFQXL \row2_buffer_reg[24][0]  ( .D(\row2_buffer[25][0] ), .CK(clk), .Q(
        \row2_buffer[24][0] ) );
  DFFQXL \row2_buffer_reg[23][0]  ( .D(\row2_buffer[24][0] ), .CK(clk), .Q(
        \row2_buffer[23][0] ) );
  DFFQXL \row2_buffer_reg[22][0]  ( .D(\row2_buffer[23][0] ), .CK(clk), .Q(
        \row2_buffer[22][0] ) );
  DFFQXL \row2_buffer_reg[21][0]  ( .D(\row2_buffer[22][0] ), .CK(clk), .Q(
        \row2_buffer[21][0] ) );
  DFFQXL \row2_buffer_reg[20][0]  ( .D(\row2_buffer[21][0] ), .CK(clk), .Q(
        \row2_buffer[20][0] ) );
  DFFQXL \row2_buffer_reg[19][0]  ( .D(\row2_buffer[20][0] ), .CK(clk), .Q(
        \row2_buffer[19][0] ) );
  DFFQXL \row2_buffer_reg[18][0]  ( .D(\row2_buffer[19][0] ), .CK(clk), .Q(
        \row2_buffer[18][0] ) );
  DFFQXL \row2_buffer_reg[17][0]  ( .D(\row2_buffer[18][0] ), .CK(clk), .Q(
        \row2_buffer[17][0] ) );
  DFFQXL \row2_buffer_reg[16][0]  ( .D(\row2_buffer[17][0] ), .CK(clk), .Q(
        \row2_buffer[16][0] ) );
  DFFQXL \row2_buffer_reg[15][0]  ( .D(\row2_buffer[16][0] ), .CK(clk), .Q(
        \row2_buffer[15][0] ) );
  DFFQXL \row2_buffer_reg[14][0]  ( .D(\row2_buffer[15][0] ), .CK(clk), .Q(
        \row2_buffer[14][0] ) );
  DFFQXL \row2_buffer_reg[13][0]  ( .D(\row2_buffer[14][0] ), .CK(clk), .Q(
        \row2_buffer[13][0] ) );
  DFFQXL \row2_buffer_reg[12][0]  ( .D(\row2_buffer[13][0] ), .CK(clk), .Q(
        \row2_buffer[12][0] ) );
  DFFQXL \row2_buffer_reg[11][0]  ( .D(\row2_buffer[12][0] ), .CK(clk), .Q(
        \row2_buffer[11][0] ) );
  DFFQXL \row2_buffer_reg[10][0]  ( .D(\row2_buffer[11][0] ), .CK(clk), .Q(
        \row2_buffer[10][0] ) );
  DFFQXL \row2_buffer_reg[9][0]  ( .D(\row2_buffer[10][0] ), .CK(clk), .Q(
        \row2_buffer[9][0] ) );
  DFFQXL \row2_buffer_reg[8][0]  ( .D(\row2_buffer[9][0] ), .CK(clk), .Q(
        \row2_buffer[8][0] ) );
  DFFQXL \row2_buffer_reg[7][0]  ( .D(\row2_buffer[8][0] ), .CK(clk), .Q(
        \row2_buffer[7][0] ) );
  DFFQXL \row2_buffer_reg[6][0]  ( .D(\row2_buffer[7][0] ), .CK(clk), .Q(
        \row2_buffer[6][0] ) );
  DFFQXL \row2_buffer_reg[5][0]  ( .D(\row2_buffer[6][0] ), .CK(clk), .Q(
        \row2_buffer[5][0] ) );
  DFFQXL \row2_buffer_reg[4][0]  ( .D(\row2_buffer[5][0] ), .CK(clk), .Q(
        \row2_buffer[4][0] ) );
  DFFQXL \row2_buffer_reg[3][0]  ( .D(\row2_buffer[4][0] ), .CK(clk), .Q(
        \row2_buffer[3][0] ) );
  DFFQXL \row1_buffer_reg[225][0]  ( .D(\row2_buffer[0][0] ), .CK(clk), .Q(
        \row1_buffer[225][0] ) );
  DFFQXL \row1_buffer_reg[224][0]  ( .D(\row1_buffer[225][0] ), .CK(clk), .Q(
        \row1_buffer[224][0] ) );
  DFFQXL \row1_buffer_reg[223][0]  ( .D(\row1_buffer[224][0] ), .CK(clk), .Q(
        \row1_buffer[223][0] ) );
  DFFQXL \row1_buffer_reg[222][0]  ( .D(\row1_buffer[223][0] ), .CK(clk), .Q(
        \row1_buffer[222][0] ) );
  DFFQXL \row1_buffer_reg[221][0]  ( .D(\row1_buffer[222][0] ), .CK(clk), .Q(
        \row1_buffer[221][0] ) );
  DFFQXL \row1_buffer_reg[220][0]  ( .D(\row1_buffer[221][0] ), .CK(clk), .Q(
        \row1_buffer[220][0] ) );
  DFFQXL \row1_buffer_reg[219][0]  ( .D(\row1_buffer[220][0] ), .CK(clk), .Q(
        \row1_buffer[219][0] ) );
  DFFQXL \row1_buffer_reg[218][0]  ( .D(\row1_buffer[219][0] ), .CK(clk), .Q(
        \row1_buffer[218][0] ) );
  DFFQXL \row1_buffer_reg[217][0]  ( .D(\row1_buffer[218][0] ), .CK(clk), .Q(
        \row1_buffer[217][0] ) );
  DFFQXL \row1_buffer_reg[216][0]  ( .D(\row1_buffer[217][0] ), .CK(clk), .Q(
        \row1_buffer[216][0] ) );
  DFFQXL \row1_buffer_reg[215][0]  ( .D(\row1_buffer[216][0] ), .CK(clk), .Q(
        \row1_buffer[215][0] ) );
  DFFQXL \row1_buffer_reg[214][0]  ( .D(\row1_buffer[215][0] ), .CK(clk), .Q(
        \row1_buffer[214][0] ) );
  DFFQXL \row1_buffer_reg[213][0]  ( .D(\row1_buffer[214][0] ), .CK(clk), .Q(
        \row1_buffer[213][0] ) );
  DFFQXL \row1_buffer_reg[212][0]  ( .D(\row1_buffer[213][0] ), .CK(clk), .Q(
        \row1_buffer[212][0] ) );
  DFFQXL \row1_buffer_reg[211][0]  ( .D(\row1_buffer[212][0] ), .CK(clk), .Q(
        \row1_buffer[211][0] ) );
  DFFQXL \row1_buffer_reg[210][0]  ( .D(\row1_buffer[211][0] ), .CK(clk), .Q(
        \row1_buffer[210][0] ) );
  DFFQXL \row1_buffer_reg[209][0]  ( .D(\row1_buffer[210][0] ), .CK(clk), .Q(
        \row1_buffer[209][0] ) );
  DFFQXL \row1_buffer_reg[208][0]  ( .D(\row1_buffer[209][0] ), .CK(clk), .Q(
        \row1_buffer[208][0] ) );
  DFFQXL \row1_buffer_reg[207][0]  ( .D(\row1_buffer[208][0] ), .CK(clk), .Q(
        \row1_buffer[207][0] ) );
  DFFQXL \row1_buffer_reg[206][0]  ( .D(\row1_buffer[207][0] ), .CK(clk), .Q(
        \row1_buffer[206][0] ) );
  DFFQXL \row1_buffer_reg[205][0]  ( .D(\row1_buffer[206][0] ), .CK(clk), .Q(
        \row1_buffer[205][0] ) );
  DFFQXL \row1_buffer_reg[204][0]  ( .D(\row1_buffer[205][0] ), .CK(clk), .Q(
        \row1_buffer[204][0] ) );
  DFFQXL \row1_buffer_reg[203][0]  ( .D(\row1_buffer[204][0] ), .CK(clk), .Q(
        \row1_buffer[203][0] ) );
  DFFQXL \row1_buffer_reg[202][0]  ( .D(\row1_buffer[203][0] ), .CK(clk), .Q(
        \row1_buffer[202][0] ) );
  DFFQXL \row1_buffer_reg[201][0]  ( .D(\row1_buffer[202][0] ), .CK(clk), .Q(
        \row1_buffer[201][0] ) );
  DFFQXL \row1_buffer_reg[200][0]  ( .D(\row1_buffer[201][0] ), .CK(clk), .Q(
        \row1_buffer[200][0] ) );
  DFFQXL \row1_buffer_reg[199][0]  ( .D(\row1_buffer[200][0] ), .CK(clk), .Q(
        \row1_buffer[199][0] ) );
  DFFQXL \row1_buffer_reg[198][0]  ( .D(\row1_buffer[199][0] ), .CK(clk), .Q(
        \row1_buffer[198][0] ) );
  DFFQXL \row1_buffer_reg[197][0]  ( .D(\row1_buffer[198][0] ), .CK(clk), .Q(
        \row1_buffer[197][0] ) );
  DFFQXL \row1_buffer_reg[196][0]  ( .D(\row1_buffer[197][0] ), .CK(clk), .Q(
        \row1_buffer[196][0] ) );
  DFFQXL \row1_buffer_reg[195][0]  ( .D(\row1_buffer[196][0] ), .CK(clk), .Q(
        \row1_buffer[195][0] ) );
  DFFQXL \row1_buffer_reg[194][0]  ( .D(\row1_buffer[195][0] ), .CK(clk), .Q(
        \row1_buffer[194][0] ) );
  DFFQXL \row1_buffer_reg[193][0]  ( .D(\row1_buffer[194][0] ), .CK(clk), .Q(
        \row1_buffer[193][0] ) );
  DFFQXL \row1_buffer_reg[192][0]  ( .D(\row1_buffer[193][0] ), .CK(clk), .Q(
        \row1_buffer[192][0] ) );
  DFFQXL \row1_buffer_reg[191][0]  ( .D(\row1_buffer[192][0] ), .CK(clk), .Q(
        \row1_buffer[191][0] ) );
  DFFQXL \row1_buffer_reg[190][0]  ( .D(\row1_buffer[191][0] ), .CK(clk), .Q(
        \row1_buffer[190][0] ) );
  DFFQXL \row1_buffer_reg[189][0]  ( .D(\row1_buffer[190][0] ), .CK(clk), .Q(
        \row1_buffer[189][0] ) );
  DFFQXL \row1_buffer_reg[188][0]  ( .D(\row1_buffer[189][0] ), .CK(clk), .Q(
        \row1_buffer[188][0] ) );
  DFFQXL \row1_buffer_reg[187][0]  ( .D(\row1_buffer[188][0] ), .CK(clk), .Q(
        \row1_buffer[187][0] ) );
  DFFQXL \row1_buffer_reg[186][0]  ( .D(\row1_buffer[187][0] ), .CK(clk), .Q(
        \row1_buffer[186][0] ) );
  DFFQXL \row1_buffer_reg[185][0]  ( .D(\row1_buffer[186][0] ), .CK(clk), .Q(
        \row1_buffer[185][0] ) );
  DFFQXL \row1_buffer_reg[184][0]  ( .D(\row1_buffer[185][0] ), .CK(clk), .Q(
        \row1_buffer[184][0] ) );
  DFFQXL \row1_buffer_reg[183][0]  ( .D(\row1_buffer[184][0] ), .CK(clk), .Q(
        \row1_buffer[183][0] ) );
  DFFQXL \row1_buffer_reg[182][0]  ( .D(\row1_buffer[183][0] ), .CK(clk), .Q(
        \row1_buffer[182][0] ) );
  DFFQXL \row1_buffer_reg[181][0]  ( .D(\row1_buffer[182][0] ), .CK(clk), .Q(
        \row1_buffer[181][0] ) );
  DFFQXL \row1_buffer_reg[180][0]  ( .D(\row1_buffer[181][0] ), .CK(clk), .Q(
        \row1_buffer[180][0] ) );
  DFFQXL \row1_buffer_reg[179][0]  ( .D(\row1_buffer[180][0] ), .CK(clk), .Q(
        \row1_buffer[179][0] ) );
  DFFQXL \row1_buffer_reg[178][0]  ( .D(\row1_buffer[179][0] ), .CK(clk), .Q(
        \row1_buffer[178][0] ) );
  DFFQXL \row1_buffer_reg[177][0]  ( .D(\row1_buffer[178][0] ), .CK(clk), .Q(
        \row1_buffer[177][0] ) );
  DFFQXL \row1_buffer_reg[176][0]  ( .D(\row1_buffer[177][0] ), .CK(clk), .Q(
        \row1_buffer[176][0] ) );
  DFFQXL \row1_buffer_reg[175][0]  ( .D(\row1_buffer[176][0] ), .CK(clk), .Q(
        \row1_buffer[175][0] ) );
  DFFQXL \row1_buffer_reg[174][0]  ( .D(\row1_buffer[175][0] ), .CK(clk), .Q(
        \row1_buffer[174][0] ) );
  DFFQXL \row1_buffer_reg[173][0]  ( .D(\row1_buffer[174][0] ), .CK(clk), .Q(
        \row1_buffer[173][0] ) );
  DFFQXL \row1_buffer_reg[172][0]  ( .D(\row1_buffer[173][0] ), .CK(clk), .Q(
        \row1_buffer[172][0] ) );
  DFFQXL \row1_buffer_reg[171][0]  ( .D(\row1_buffer[172][0] ), .CK(clk), .Q(
        \row1_buffer[171][0] ) );
  DFFQXL \row1_buffer_reg[170][0]  ( .D(\row1_buffer[171][0] ), .CK(clk), .Q(
        \row1_buffer[170][0] ) );
  DFFQXL \row1_buffer_reg[169][0]  ( .D(\row1_buffer[170][0] ), .CK(clk), .Q(
        \row1_buffer[169][0] ) );
  DFFQXL \row1_buffer_reg[168][0]  ( .D(\row1_buffer[169][0] ), .CK(clk), .Q(
        \row1_buffer[168][0] ) );
  DFFQXL \row1_buffer_reg[167][0]  ( .D(\row1_buffer[168][0] ), .CK(clk), .Q(
        \row1_buffer[167][0] ) );
  DFFQXL \row1_buffer_reg[166][0]  ( .D(\row1_buffer[167][0] ), .CK(clk), .Q(
        \row1_buffer[166][0] ) );
  DFFQXL \row1_buffer_reg[165][0]  ( .D(\row1_buffer[166][0] ), .CK(clk), .Q(
        \row1_buffer[165][0] ) );
  DFFQXL \row1_buffer_reg[164][0]  ( .D(\row1_buffer[165][0] ), .CK(clk), .Q(
        \row1_buffer[164][0] ) );
  DFFQXL \row1_buffer_reg[163][0]  ( .D(\row1_buffer[164][0] ), .CK(clk), .Q(
        \row1_buffer[163][0] ) );
  DFFQXL \row1_buffer_reg[162][0]  ( .D(\row1_buffer[163][0] ), .CK(clk), .Q(
        \row1_buffer[162][0] ) );
  DFFQXL \row1_buffer_reg[161][0]  ( .D(\row1_buffer[162][0] ), .CK(clk), .Q(
        \row1_buffer[161][0] ) );
  DFFQXL \row1_buffer_reg[160][0]  ( .D(\row1_buffer[161][0] ), .CK(clk), .Q(
        \row1_buffer[160][0] ) );
  DFFQXL \row1_buffer_reg[159][0]  ( .D(\row1_buffer[160][0] ), .CK(clk), .Q(
        \row1_buffer[159][0] ) );
  DFFQXL \row1_buffer_reg[158][0]  ( .D(\row1_buffer[159][0] ), .CK(clk), .Q(
        \row1_buffer[158][0] ) );
  DFFQXL \row1_buffer_reg[157][0]  ( .D(\row1_buffer[158][0] ), .CK(clk), .Q(
        \row1_buffer[157][0] ) );
  DFFQXL \row1_buffer_reg[156][0]  ( .D(\row1_buffer[157][0] ), .CK(clk), .Q(
        \row1_buffer[156][0] ) );
  DFFQXL \row1_buffer_reg[155][0]  ( .D(\row1_buffer[156][0] ), .CK(clk), .Q(
        \row1_buffer[155][0] ) );
  DFFQXL \row1_buffer_reg[154][0]  ( .D(\row1_buffer[155][0] ), .CK(clk), .Q(
        \row1_buffer[154][0] ) );
  DFFQXL \row1_buffer_reg[153][0]  ( .D(\row1_buffer[154][0] ), .CK(clk), .Q(
        \row1_buffer[153][0] ) );
  DFFQXL \row1_buffer_reg[152][0]  ( .D(\row1_buffer[153][0] ), .CK(clk), .Q(
        \row1_buffer[152][0] ) );
  DFFQXL \row1_buffer_reg[151][0]  ( .D(\row1_buffer[152][0] ), .CK(clk), .Q(
        \row1_buffer[151][0] ) );
  DFFQXL \row1_buffer_reg[150][0]  ( .D(\row1_buffer[151][0] ), .CK(clk), .Q(
        \row1_buffer[150][0] ) );
  DFFQXL \row1_buffer_reg[149][0]  ( .D(\row1_buffer[150][0] ), .CK(clk), .Q(
        \row1_buffer[149][0] ) );
  DFFQXL \row1_buffer_reg[148][0]  ( .D(\row1_buffer[149][0] ), .CK(clk), .Q(
        \row1_buffer[148][0] ) );
  DFFQXL \row1_buffer_reg[147][0]  ( .D(\row1_buffer[148][0] ), .CK(clk), .Q(
        \row1_buffer[147][0] ) );
  DFFQXL \row1_buffer_reg[146][0]  ( .D(\row1_buffer[147][0] ), .CK(clk), .Q(
        \row1_buffer[146][0] ) );
  DFFQXL \row1_buffer_reg[145][0]  ( .D(\row1_buffer[146][0] ), .CK(clk), .Q(
        \row1_buffer[145][0] ) );
  DFFQXL \row1_buffer_reg[144][0]  ( .D(\row1_buffer[145][0] ), .CK(clk), .Q(
        \row1_buffer[144][0] ) );
  DFFQXL \row1_buffer_reg[143][0]  ( .D(\row1_buffer[144][0] ), .CK(clk), .Q(
        \row1_buffer[143][0] ) );
  DFFQXL \row1_buffer_reg[142][0]  ( .D(\row1_buffer[143][0] ), .CK(clk), .Q(
        \row1_buffer[142][0] ) );
  DFFQXL \row1_buffer_reg[141][0]  ( .D(\row1_buffer[142][0] ), .CK(clk), .Q(
        \row1_buffer[141][0] ) );
  DFFQXL \row1_buffer_reg[140][0]  ( .D(\row1_buffer[141][0] ), .CK(clk), .Q(
        \row1_buffer[140][0] ) );
  DFFQXL \row1_buffer_reg[139][0]  ( .D(\row1_buffer[140][0] ), .CK(clk), .Q(
        \row1_buffer[139][0] ) );
  DFFQXL \row1_buffer_reg[138][0]  ( .D(\row1_buffer[139][0] ), .CK(clk), .Q(
        \row1_buffer[138][0] ) );
  DFFQXL \row1_buffer_reg[137][0]  ( .D(\row1_buffer[138][0] ), .CK(clk), .Q(
        \row1_buffer[137][0] ) );
  DFFQXL \row1_buffer_reg[136][0]  ( .D(\row1_buffer[137][0] ), .CK(clk), .Q(
        \row1_buffer[136][0] ) );
  DFFQXL \row1_buffer_reg[135][0]  ( .D(\row1_buffer[136][0] ), .CK(clk), .Q(
        \row1_buffer[135][0] ) );
  DFFQXL \row1_buffer_reg[134][0]  ( .D(\row1_buffer[135][0] ), .CK(clk), .Q(
        \row1_buffer[134][0] ) );
  DFFQXL \row1_buffer_reg[133][0]  ( .D(\row1_buffer[134][0] ), .CK(clk), .Q(
        \row1_buffer[133][0] ) );
  DFFQXL \row1_buffer_reg[132][0]  ( .D(\row1_buffer[133][0] ), .CK(clk), .Q(
        \row1_buffer[132][0] ) );
  DFFQXL \row1_buffer_reg[131][0]  ( .D(\row1_buffer[132][0] ), .CK(clk), .Q(
        \row1_buffer[131][0] ) );
  DFFQXL \row1_buffer_reg[130][0]  ( .D(\row1_buffer[131][0] ), .CK(clk), .Q(
        \row1_buffer[130][0] ) );
  DFFQXL \row1_buffer_reg[129][0]  ( .D(\row1_buffer[130][0] ), .CK(clk), .Q(
        \row1_buffer[129][0] ) );
  DFFQXL \row1_buffer_reg[128][0]  ( .D(\row1_buffer[129][0] ), .CK(clk), .Q(
        \row1_buffer[128][0] ) );
  DFFQXL \row1_buffer_reg[127][0]  ( .D(\row1_buffer[128][0] ), .CK(clk), .Q(
        \row1_buffer[127][0] ) );
  DFFQXL \row1_buffer_reg[126][0]  ( .D(\row1_buffer[127][0] ), .CK(clk), .Q(
        \row1_buffer[126][0] ) );
  DFFQXL \row1_buffer_reg[125][0]  ( .D(\row1_buffer[126][0] ), .CK(clk), .Q(
        \row1_buffer[125][0] ) );
  DFFQXL \row1_buffer_reg[124][0]  ( .D(\row1_buffer[125][0] ), .CK(clk), .Q(
        \row1_buffer[124][0] ) );
  DFFQXL \row1_buffer_reg[123][0]  ( .D(\row1_buffer[124][0] ), .CK(clk), .Q(
        \row1_buffer[123][0] ) );
  DFFQXL \row1_buffer_reg[122][0]  ( .D(\row1_buffer[123][0] ), .CK(clk), .Q(
        \row1_buffer[122][0] ) );
  DFFQXL \row1_buffer_reg[121][0]  ( .D(\row1_buffer[122][0] ), .CK(clk), .Q(
        \row1_buffer[121][0] ) );
  DFFQXL \row1_buffer_reg[120][0]  ( .D(\row1_buffer[121][0] ), .CK(clk), .Q(
        \row1_buffer[120][0] ) );
  DFFQXL \row1_buffer_reg[119][0]  ( .D(\row1_buffer[120][0] ), .CK(clk), .Q(
        \row1_buffer[119][0] ) );
  DFFQXL \row1_buffer_reg[118][0]  ( .D(\row1_buffer[119][0] ), .CK(clk), .Q(
        \row1_buffer[118][0] ) );
  DFFQXL \row1_buffer_reg[117][0]  ( .D(\row1_buffer[118][0] ), .CK(clk), .Q(
        \row1_buffer[117][0] ) );
  DFFQXL \row1_buffer_reg[116][0]  ( .D(\row1_buffer[117][0] ), .CK(clk), .Q(
        \row1_buffer[116][0] ) );
  DFFQXL \row1_buffer_reg[115][0]  ( .D(\row1_buffer[116][0] ), .CK(clk), .Q(
        \row1_buffer[115][0] ) );
  DFFQXL \row1_buffer_reg[114][0]  ( .D(\row1_buffer[115][0] ), .CK(clk), .Q(
        \row1_buffer[114][0] ) );
  DFFQXL \row1_buffer_reg[113][0]  ( .D(\row1_buffer[114][0] ), .CK(clk), .Q(
        \row1_buffer[113][0] ) );
  DFFQXL \row1_buffer_reg[112][0]  ( .D(\row1_buffer[113][0] ), .CK(clk), .Q(
        \row1_buffer[112][0] ) );
  DFFQXL \row1_buffer_reg[111][0]  ( .D(\row1_buffer[112][0] ), .CK(clk), .Q(
        \row1_buffer[111][0] ) );
  DFFQXL \row1_buffer_reg[110][0]  ( .D(\row1_buffer[111][0] ), .CK(clk), .Q(
        \row1_buffer[110][0] ) );
  DFFQXL \row1_buffer_reg[109][0]  ( .D(\row1_buffer[110][0] ), .CK(clk), .Q(
        \row1_buffer[109][0] ) );
  DFFQXL \row1_buffer_reg[108][0]  ( .D(\row1_buffer[109][0] ), .CK(clk), .Q(
        \row1_buffer[108][0] ) );
  DFFQXL \row1_buffer_reg[107][0]  ( .D(\row1_buffer[108][0] ), .CK(clk), .Q(
        \row1_buffer[107][0] ) );
  DFFQXL \row1_buffer_reg[106][0]  ( .D(\row1_buffer[107][0] ), .CK(clk), .Q(
        \row1_buffer[106][0] ) );
  DFFQXL \row1_buffer_reg[105][0]  ( .D(\row1_buffer[106][0] ), .CK(clk), .Q(
        \row1_buffer[105][0] ) );
  DFFQXL \row1_buffer_reg[104][0]  ( .D(\row1_buffer[105][0] ), .CK(clk), .Q(
        \row1_buffer[104][0] ) );
  DFFQXL \row1_buffer_reg[103][0]  ( .D(\row1_buffer[104][0] ), .CK(clk), .Q(
        \row1_buffer[103][0] ) );
  DFFQXL \row1_buffer_reg[102][0]  ( .D(\row1_buffer[103][0] ), .CK(clk), .Q(
        \row1_buffer[102][0] ) );
  DFFQXL \row1_buffer_reg[101][0]  ( .D(\row1_buffer[102][0] ), .CK(clk), .Q(
        \row1_buffer[101][0] ) );
  DFFQXL \row1_buffer_reg[100][0]  ( .D(\row1_buffer[101][0] ), .CK(clk), .Q(
        \row1_buffer[100][0] ) );
  DFFQXL \row1_buffer_reg[99][0]  ( .D(\row1_buffer[100][0] ), .CK(clk), .Q(
        \row1_buffer[99][0] ) );
  DFFQXL \row1_buffer_reg[98][0]  ( .D(\row1_buffer[99][0] ), .CK(clk), .Q(
        \row1_buffer[98][0] ) );
  DFFQXL \row1_buffer_reg[97][0]  ( .D(\row1_buffer[98][0] ), .CK(clk), .Q(
        \row1_buffer[97][0] ) );
  DFFQXL \row1_buffer_reg[96][0]  ( .D(\row1_buffer[97][0] ), .CK(clk), .Q(
        \row1_buffer[96][0] ) );
  DFFQXL \row1_buffer_reg[95][0]  ( .D(\row1_buffer[96][0] ), .CK(clk), .Q(
        \row1_buffer[95][0] ) );
  DFFQXL \row1_buffer_reg[94][0]  ( .D(\row1_buffer[95][0] ), .CK(clk), .Q(
        \row1_buffer[94][0] ) );
  DFFQXL \row1_buffer_reg[93][0]  ( .D(\row1_buffer[94][0] ), .CK(clk), .Q(
        \row1_buffer[93][0] ) );
  DFFQXL \row1_buffer_reg[92][0]  ( .D(\row1_buffer[93][0] ), .CK(clk), .Q(
        \row1_buffer[92][0] ) );
  DFFQXL \row1_buffer_reg[91][0]  ( .D(\row1_buffer[92][0] ), .CK(clk), .Q(
        \row1_buffer[91][0] ) );
  DFFQXL \row1_buffer_reg[90][0]  ( .D(\row1_buffer[91][0] ), .CK(clk), .Q(
        \row1_buffer[90][0] ) );
  DFFQXL \row1_buffer_reg[89][0]  ( .D(\row1_buffer[90][0] ), .CK(clk), .Q(
        \row1_buffer[89][0] ) );
  DFFQXL \row1_buffer_reg[88][0]  ( .D(\row1_buffer[89][0] ), .CK(clk), .Q(
        \row1_buffer[88][0] ) );
  DFFQXL \row1_buffer_reg[87][0]  ( .D(\row1_buffer[88][0] ), .CK(clk), .Q(
        \row1_buffer[87][0] ) );
  DFFQXL \row1_buffer_reg[86][0]  ( .D(\row1_buffer[87][0] ), .CK(clk), .Q(
        \row1_buffer[86][0] ) );
  DFFQXL \row1_buffer_reg[85][0]  ( .D(\row1_buffer[86][0] ), .CK(clk), .Q(
        \row1_buffer[85][0] ) );
  DFFQXL \row1_buffer_reg[84][0]  ( .D(\row1_buffer[85][0] ), .CK(clk), .Q(
        \row1_buffer[84][0] ) );
  DFFQXL \row1_buffer_reg[83][0]  ( .D(\row1_buffer[84][0] ), .CK(clk), .Q(
        \row1_buffer[83][0] ) );
  DFFQXL \row1_buffer_reg[82][0]  ( .D(\row1_buffer[83][0] ), .CK(clk), .Q(
        \row1_buffer[82][0] ) );
  DFFQXL \row1_buffer_reg[81][0]  ( .D(\row1_buffer[82][0] ), .CK(clk), .Q(
        \row1_buffer[81][0] ) );
  DFFQXL \row1_buffer_reg[80][0]  ( .D(\row1_buffer[81][0] ), .CK(clk), .Q(
        \row1_buffer[80][0] ) );
  DFFQXL \row1_buffer_reg[79][0]  ( .D(\row1_buffer[80][0] ), .CK(clk), .Q(
        \row1_buffer[79][0] ) );
  DFFQXL \row1_buffer_reg[78][0]  ( .D(\row1_buffer[79][0] ), .CK(clk), .Q(
        \row1_buffer[78][0] ) );
  DFFQXL \row1_buffer_reg[77][0]  ( .D(\row1_buffer[78][0] ), .CK(clk), .Q(
        \row1_buffer[77][0] ) );
  DFFQXL \row1_buffer_reg[76][0]  ( .D(\row1_buffer[77][0] ), .CK(clk), .Q(
        \row1_buffer[76][0] ) );
  DFFQXL \row1_buffer_reg[75][0]  ( .D(\row1_buffer[76][0] ), .CK(clk), .Q(
        \row1_buffer[75][0] ) );
  DFFQXL \row1_buffer_reg[74][0]  ( .D(\row1_buffer[75][0] ), .CK(clk), .Q(
        \row1_buffer[74][0] ) );
  DFFQXL \row1_buffer_reg[73][0]  ( .D(\row1_buffer[74][0] ), .CK(clk), .Q(
        \row1_buffer[73][0] ) );
  DFFQXL \row1_buffer_reg[72][0]  ( .D(\row1_buffer[73][0] ), .CK(clk), .Q(
        \row1_buffer[72][0] ) );
  DFFQXL \row1_buffer_reg[71][0]  ( .D(\row1_buffer[72][0] ), .CK(clk), .Q(
        \row1_buffer[71][0] ) );
  DFFQXL \row1_buffer_reg[70][0]  ( .D(\row1_buffer[71][0] ), .CK(clk), .Q(
        \row1_buffer[70][0] ) );
  DFFQXL \row1_buffer_reg[69][0]  ( .D(\row1_buffer[70][0] ), .CK(clk), .Q(
        \row1_buffer[69][0] ) );
  DFFQXL \row1_buffer_reg[68][0]  ( .D(\row1_buffer[69][0] ), .CK(clk), .Q(
        \row1_buffer[68][0] ) );
  DFFQXL \row1_buffer_reg[67][0]  ( .D(\row1_buffer[68][0] ), .CK(clk), .Q(
        \row1_buffer[67][0] ) );
  DFFQXL \row1_buffer_reg[66][0]  ( .D(\row1_buffer[67][0] ), .CK(clk), .Q(
        \row1_buffer[66][0] ) );
  DFFQXL \row1_buffer_reg[65][0]  ( .D(\row1_buffer[66][0] ), .CK(clk), .Q(
        \row1_buffer[65][0] ) );
  DFFQXL \row1_buffer_reg[64][0]  ( .D(\row1_buffer[65][0] ), .CK(clk), .Q(
        \row1_buffer[64][0] ) );
  DFFQXL \row1_buffer_reg[63][0]  ( .D(\row1_buffer[64][0] ), .CK(clk), .Q(
        \row1_buffer[63][0] ) );
  DFFQXL \row1_buffer_reg[62][0]  ( .D(\row1_buffer[63][0] ), .CK(clk), .Q(
        \row1_buffer[62][0] ) );
  DFFQXL \row1_buffer_reg[61][0]  ( .D(\row1_buffer[62][0] ), .CK(clk), .Q(
        \row1_buffer[61][0] ) );
  DFFQXL \row1_buffer_reg[60][0]  ( .D(\row1_buffer[61][0] ), .CK(clk), .Q(
        \row1_buffer[60][0] ) );
  DFFQXL \row1_buffer_reg[59][0]  ( .D(\row1_buffer[60][0] ), .CK(clk), .Q(
        \row1_buffer[59][0] ) );
  DFFQXL \row1_buffer_reg[58][0]  ( .D(\row1_buffer[59][0] ), .CK(clk), .Q(
        \row1_buffer[58][0] ) );
  DFFQXL \row1_buffer_reg[57][0]  ( .D(\row1_buffer[58][0] ), .CK(clk), .Q(
        \row1_buffer[57][0] ) );
  DFFQXL \row1_buffer_reg[56][0]  ( .D(\row1_buffer[57][0] ), .CK(clk), .Q(
        \row1_buffer[56][0] ) );
  DFFQXL \row1_buffer_reg[55][0]  ( .D(\row1_buffer[56][0] ), .CK(clk), .Q(
        \row1_buffer[55][0] ) );
  DFFQXL \row1_buffer_reg[54][0]  ( .D(\row1_buffer[55][0] ), .CK(clk), .Q(
        \row1_buffer[54][0] ) );
  DFFQXL \row1_buffer_reg[53][0]  ( .D(\row1_buffer[54][0] ), .CK(clk), .Q(
        \row1_buffer[53][0] ) );
  DFFQXL \row1_buffer_reg[52][0]  ( .D(\row1_buffer[53][0] ), .CK(clk), .Q(
        \row1_buffer[52][0] ) );
  DFFQXL \row1_buffer_reg[51][0]  ( .D(\row1_buffer[52][0] ), .CK(clk), .Q(
        \row1_buffer[51][0] ) );
  DFFQXL \row1_buffer_reg[50][0]  ( .D(\row1_buffer[51][0] ), .CK(clk), .Q(
        \row1_buffer[50][0] ) );
  DFFQXL \row1_buffer_reg[49][0]  ( .D(\row1_buffer[50][0] ), .CK(clk), .Q(
        \row1_buffer[49][0] ) );
  DFFQXL \row1_buffer_reg[48][0]  ( .D(\row1_buffer[49][0] ), .CK(clk), .Q(
        \row1_buffer[48][0] ) );
  DFFQXL \row1_buffer_reg[47][0]  ( .D(\row1_buffer[48][0] ), .CK(clk), .Q(
        \row1_buffer[47][0] ) );
  DFFQXL \row1_buffer_reg[46][0]  ( .D(\row1_buffer[47][0] ), .CK(clk), .Q(
        \row1_buffer[46][0] ) );
  DFFQXL \row1_buffer_reg[45][0]  ( .D(\row1_buffer[46][0] ), .CK(clk), .Q(
        \row1_buffer[45][0] ) );
  DFFQXL \row1_buffer_reg[44][0]  ( .D(\row1_buffer[45][0] ), .CK(clk), .Q(
        \row1_buffer[44][0] ) );
  DFFQXL \row1_buffer_reg[43][0]  ( .D(\row1_buffer[44][0] ), .CK(clk), .Q(
        \row1_buffer[43][0] ) );
  DFFQXL \row1_buffer_reg[42][0]  ( .D(\row1_buffer[43][0] ), .CK(clk), .Q(
        \row1_buffer[42][0] ) );
  DFFQXL \row1_buffer_reg[41][0]  ( .D(\row1_buffer[42][0] ), .CK(clk), .Q(
        \row1_buffer[41][0] ) );
  DFFQXL \row1_buffer_reg[40][0]  ( .D(\row1_buffer[41][0] ), .CK(clk), .Q(
        \row1_buffer[40][0] ) );
  DFFQXL \row1_buffer_reg[39][0]  ( .D(\row1_buffer[40][0] ), .CK(clk), .Q(
        \row1_buffer[39][0] ) );
  DFFQXL \row1_buffer_reg[38][0]  ( .D(\row1_buffer[39][0] ), .CK(clk), .Q(
        \row1_buffer[38][0] ) );
  DFFQXL \row1_buffer_reg[37][0]  ( .D(\row1_buffer[38][0] ), .CK(clk), .Q(
        \row1_buffer[37][0] ) );
  DFFQXL \row1_buffer_reg[36][0]  ( .D(\row1_buffer[37][0] ), .CK(clk), .Q(
        \row1_buffer[36][0] ) );
  DFFQXL \row1_buffer_reg[35][0]  ( .D(\row1_buffer[36][0] ), .CK(clk), .Q(
        \row1_buffer[35][0] ) );
  DFFQXL \row1_buffer_reg[34][0]  ( .D(\row1_buffer[35][0] ), .CK(clk), .Q(
        \row1_buffer[34][0] ) );
  DFFQXL \row1_buffer_reg[33][0]  ( .D(\row1_buffer[34][0] ), .CK(clk), .Q(
        \row1_buffer[33][0] ) );
  DFFQXL \row1_buffer_reg[32][0]  ( .D(\row1_buffer[33][0] ), .CK(clk), .Q(
        \row1_buffer[32][0] ) );
  DFFQXL \row1_buffer_reg[31][0]  ( .D(\row1_buffer[32][0] ), .CK(clk), .Q(
        \row1_buffer[31][0] ) );
  DFFQXL \row1_buffer_reg[30][0]  ( .D(\row1_buffer[31][0] ), .CK(clk), .Q(
        \row1_buffer[30][0] ) );
  DFFQXL \row1_buffer_reg[29][0]  ( .D(\row1_buffer[30][0] ), .CK(clk), .Q(
        \row1_buffer[29][0] ) );
  DFFQXL \row1_buffer_reg[28][0]  ( .D(\row1_buffer[29][0] ), .CK(clk), .Q(
        \row1_buffer[28][0] ) );
  DFFQXL \row1_buffer_reg[27][0]  ( .D(\row1_buffer[28][0] ), .CK(clk), .Q(
        \row1_buffer[27][0] ) );
  DFFQXL \row1_buffer_reg[26][0]  ( .D(\row1_buffer[27][0] ), .CK(clk), .Q(
        \row1_buffer[26][0] ) );
  DFFQXL \row1_buffer_reg[25][0]  ( .D(\row1_buffer[26][0] ), .CK(clk), .Q(
        \row1_buffer[25][0] ) );
  DFFQXL \row1_buffer_reg[24][0]  ( .D(\row1_buffer[25][0] ), .CK(clk), .Q(
        \row1_buffer[24][0] ) );
  DFFQXL \row1_buffer_reg[23][0]  ( .D(\row1_buffer[24][0] ), .CK(clk), .Q(
        \row1_buffer[23][0] ) );
  DFFQXL \row1_buffer_reg[22][0]  ( .D(\row1_buffer[23][0] ), .CK(clk), .Q(
        \row1_buffer[22][0] ) );
  DFFQXL \row1_buffer_reg[21][0]  ( .D(\row1_buffer[22][0] ), .CK(clk), .Q(
        \row1_buffer[21][0] ) );
  DFFQXL \row1_buffer_reg[20][0]  ( .D(\row1_buffer[21][0] ), .CK(clk), .Q(
        \row1_buffer[20][0] ) );
  DFFQXL \row1_buffer_reg[19][0]  ( .D(\row1_buffer[20][0] ), .CK(clk), .Q(
        \row1_buffer[19][0] ) );
  DFFQXL \row1_buffer_reg[18][0]  ( .D(\row1_buffer[19][0] ), .CK(clk), .Q(
        \row1_buffer[18][0] ) );
  DFFQXL \row1_buffer_reg[17][0]  ( .D(\row1_buffer[18][0] ), .CK(clk), .Q(
        \row1_buffer[17][0] ) );
  DFFQXL \row1_buffer_reg[16][0]  ( .D(\row1_buffer[17][0] ), .CK(clk), .Q(
        \row1_buffer[16][0] ) );
  DFFQXL \row1_buffer_reg[15][0]  ( .D(\row1_buffer[16][0] ), .CK(clk), .Q(
        \row1_buffer[15][0] ) );
  DFFQXL \row1_buffer_reg[14][0]  ( .D(\row1_buffer[15][0] ), .CK(clk), .Q(
        \row1_buffer[14][0] ) );
  DFFQXL \row1_buffer_reg[13][0]  ( .D(\row1_buffer[14][0] ), .CK(clk), .Q(
        \row1_buffer[13][0] ) );
  DFFQXL \row1_buffer_reg[12][0]  ( .D(\row1_buffer[13][0] ), .CK(clk), .Q(
        \row1_buffer[12][0] ) );
  DFFQXL \row1_buffer_reg[11][0]  ( .D(\row1_buffer[12][0] ), .CK(clk), .Q(
        \row1_buffer[11][0] ) );
  DFFQXL \row1_buffer_reg[10][0]  ( .D(\row1_buffer[11][0] ), .CK(clk), .Q(
        \row1_buffer[10][0] ) );
  DFFQXL \row1_buffer_reg[9][0]  ( .D(\row1_buffer[10][0] ), .CK(clk), .Q(
        \row1_buffer[9][0] ) );
  DFFQXL \row1_buffer_reg[8][0]  ( .D(\row1_buffer[9][0] ), .CK(clk), .Q(
        \row1_buffer[8][0] ) );
  DFFQXL \row1_buffer_reg[7][0]  ( .D(\row1_buffer[8][0] ), .CK(clk), .Q(
        \row1_buffer[7][0] ) );
  DFFQXL \row1_buffer_reg[6][0]  ( .D(\row1_buffer[7][0] ), .CK(clk), .Q(
        \row1_buffer[6][0] ) );
  DFFQXL \row1_buffer_reg[5][0]  ( .D(\row1_buffer[6][0] ), .CK(clk), .Q(
        \row1_buffer[5][0] ) );
  DFFQXL \row1_buffer_reg[4][0]  ( .D(\row1_buffer[5][0] ), .CK(clk), .Q(
        \row1_buffer[4][0] ) );
  DFFQXL \row1_buffer_reg[3][0]  ( .D(\row1_buffer[4][0] ), .CK(clk), .Q(
        \row1_buffer[3][0] ) );
  DFFQXL \row3_buffer_reg[2][6]  ( .D(in_pixel[6]), .CK(clk), .Q(
        \row3_buffer[2][6] ) );
  DFFQXL \row3_buffer_reg[1][6]  ( .D(\row3_buffer[2][6] ), .CK(clk), .Q(
        \row3_buffer[1][6] ) );
  DFFQXL \row3_buffer_reg[0][6]  ( .D(\row3_buffer[1][6] ), .CK(clk), .Q(
        \row3_buffer[0][6] ) );
  DFFQXL \row2_buffer_reg[2][6]  ( .D(\row2_buffer[3][6] ), .CK(clk), .Q(
        \row2_buffer[2][6] ) );
  DFFQXL \row2_buffer_reg[1][6]  ( .D(\row2_buffer[2][6] ), .CK(clk), .Q(
        \row2_buffer[1][6] ) );
  DFFQXL \row2_buffer_reg[0][6]  ( .D(\row2_buffer[1][6] ), .CK(clk), .Q(
        \row2_buffer[0][6] ) );
  DFFQXL \row1_buffer_reg[2][6]  ( .D(\row1_buffer[3][6] ), .CK(clk), .Q(
        \row1_buffer[2][6] ) );
  DFFQXL \row1_buffer_reg[1][6]  ( .D(\row1_buffer[2][6] ), .CK(clk), .Q(
        \row1_buffer[1][6] ) );
  DFFQXL \row3_buffer_reg[2][4]  ( .D(in_pixel[4]), .CK(clk), .Q(
        \row3_buffer[2][4] ) );
  DFFQXL \row3_buffer_reg[1][4]  ( .D(\row3_buffer[2][4] ), .CK(clk), .Q(
        \row3_buffer[1][4] ) );
  DFFQXL \row3_buffer_reg[0][4]  ( .D(\row3_buffer[1][4] ), .CK(clk), .Q(
        \row3_buffer[0][4] ) );
  DFFQXL \row2_buffer_reg[2][4]  ( .D(\row2_buffer[3][4] ), .CK(clk), .Q(
        \row2_buffer[2][4] ) );
  DFFQXL \row2_buffer_reg[1][4]  ( .D(\row2_buffer[2][4] ), .CK(clk), .Q(
        \row2_buffer[1][4] ) );
  DFFQXL \row2_buffer_reg[0][4]  ( .D(\row2_buffer[1][4] ), .CK(clk), .Q(
        \row2_buffer[0][4] ) );
  DFFQXL \row1_buffer_reg[2][4]  ( .D(\row1_buffer[3][4] ), .CK(clk), .Q(
        \row1_buffer[2][4] ) );
  DFFQXL \row1_buffer_reg[1][4]  ( .D(\row1_buffer[2][4] ), .CK(clk), .Q(
        \row1_buffer[1][4] ) );
  DFFQXL \row3_buffer_reg[2][2]  ( .D(in_pixel[2]), .CK(clk), .Q(
        \row3_buffer[2][2] ) );
  DFFQXL \row3_buffer_reg[1][2]  ( .D(\row3_buffer[2][2] ), .CK(clk), .Q(
        \row3_buffer[1][2] ) );
  DFFQXL \row3_buffer_reg[0][2]  ( .D(\row3_buffer[1][2] ), .CK(clk), .Q(
        \row3_buffer[0][2] ) );
  DFFQXL \row2_buffer_reg[2][2]  ( .D(\row2_buffer[3][2] ), .CK(clk), .Q(
        \row2_buffer[2][2] ) );
  DFFQXL \row2_buffer_reg[1][2]  ( .D(\row2_buffer[2][2] ), .CK(clk), .Q(
        \row2_buffer[1][2] ) );
  DFFQXL \row2_buffer_reg[0][2]  ( .D(\row2_buffer[1][2] ), .CK(clk), .Q(
        \row2_buffer[0][2] ) );
  DFFQXL \row1_buffer_reg[2][2]  ( .D(\row1_buffer[3][2] ), .CK(clk), .Q(
        \row1_buffer[2][2] ) );
  DFFQXL \row1_buffer_reg[1][2]  ( .D(\row1_buffer[2][2] ), .CK(clk), .Q(
        \row1_buffer[1][2] ) );
  DFFQXL \row3_buffer_reg[2][1]  ( .D(in_pixel[1]), .CK(clk), .Q(
        \row3_buffer[2][1] ) );
  DFFQXL \row3_buffer_reg[1][1]  ( .D(\row3_buffer[2][1] ), .CK(clk), .Q(
        \row3_buffer[1][1] ) );
  DFFQXL \row3_buffer_reg[0][1]  ( .D(\row3_buffer[1][1] ), .CK(clk), .Q(
        \row3_buffer[0][1] ) );
  DFFQXL \row2_buffer_reg[2][1]  ( .D(\row2_buffer[3][1] ), .CK(clk), .Q(
        \row2_buffer[2][1] ) );
  DFFQXL \row2_buffer_reg[1][1]  ( .D(\row2_buffer[2][1] ), .CK(clk), .Q(
        \row2_buffer[1][1] ) );
  DFFQXL \row2_buffer_reg[0][1]  ( .D(\row2_buffer[1][1] ), .CK(clk), .Q(
        \row2_buffer[0][1] ) );
  DFFQXL \row1_buffer_reg[2][1]  ( .D(\row1_buffer[3][1] ), .CK(clk), .Q(
        \row1_buffer[2][1] ) );
  DFFQXL \row1_buffer_reg[1][1]  ( .D(\row1_buffer[2][1] ), .CK(clk), .Q(
        \row1_buffer[1][1] ) );
  DFFQXL \row3_buffer_reg[2][0]  ( .D(in_pixel[0]), .CK(clk), .Q(
        \row3_buffer[2][0] ) );
  DFFQXL \row3_buffer_reg[1][0]  ( .D(\row3_buffer[2][0] ), .CK(clk), .Q(
        \row3_buffer[1][0] ) );
  DFFQXL \row3_buffer_reg[0][0]  ( .D(\row3_buffer[1][0] ), .CK(clk), .Q(
        \row3_buffer[0][0] ) );
  DFFQXL \row2_buffer_reg[2][0]  ( .D(\row2_buffer[3][0] ), .CK(clk), .Q(
        \row2_buffer[2][0] ) );
  DFFQXL \row2_buffer_reg[1][0]  ( .D(\row2_buffer[2][0] ), .CK(clk), .Q(
        \row2_buffer[1][0] ) );
  DFFQXL \row2_buffer_reg[0][0]  ( .D(\row2_buffer[1][0] ), .CK(clk), .Q(
        \row2_buffer[0][0] ) );
  DFFQXL \row1_buffer_reg[2][0]  ( .D(\row1_buffer[3][0] ), .CK(clk), .Q(
        \row1_buffer[2][0] ) );
  DFFQXL \row1_buffer_reg[1][0]  ( .D(\row1_buffer[2][0] ), .CK(clk), .Q(
        \row1_buffer[1][0] ) );
  DFFQXL \row3_buffer_reg[2][7]  ( .D(in_pixel[7]), .CK(clk), .Q(
        \row3_buffer[2][7] ) );
  DFFQXL \row3_buffer_reg[1][7]  ( .D(\row3_buffer[2][7] ), .CK(clk), .Q(
        \row3_buffer[1][7] ) );
  DFFQXL \row3_buffer_reg[0][7]  ( .D(\row3_buffer[1][7] ), .CK(clk), .Q(
        \row3_buffer[0][7] ) );
  DFFQXL \row2_buffer_reg[2][7]  ( .D(\row2_buffer[3][7] ), .CK(clk), .Q(
        \row2_buffer[2][7] ) );
  DFFQXL \row2_buffer_reg[1][7]  ( .D(\row2_buffer[2][7] ), .CK(clk), .Q(
        \row2_buffer[1][7] ) );
  DFFQXL \row2_buffer_reg[0][7]  ( .D(\row2_buffer[1][7] ), .CK(clk), .Q(
        \row2_buffer[0][7] ) );
  DFFQXL \row1_buffer_reg[2][7]  ( .D(\row1_buffer[3][7] ), .CK(clk), .Q(
        \row1_buffer[2][7] ) );
  DFFQXL \row1_buffer_reg[1][7]  ( .D(\row1_buffer[2][7] ), .CK(clk), .Q(
        \row1_buffer[1][7] ) );
  DFFQXL \row3_buffer_reg[2][5]  ( .D(in_pixel[5]), .CK(clk), .Q(
        \row3_buffer[2][5] ) );
  DFFQXL \row3_buffer_reg[1][5]  ( .D(\row3_buffer[2][5] ), .CK(clk), .Q(
        \row3_buffer[1][5] ) );
  DFFQXL \row3_buffer_reg[0][5]  ( .D(\row3_buffer[1][5] ), .CK(clk), .Q(
        \row3_buffer[0][5] ) );
  DFFQXL \row2_buffer_reg[2][5]  ( .D(\row2_buffer[3][5] ), .CK(clk), .Q(
        \row2_buffer[2][5] ) );
  DFFQXL \row2_buffer_reg[1][5]  ( .D(\row2_buffer[2][5] ), .CK(clk), .Q(
        \row2_buffer[1][5] ) );
  DFFQXL \row2_buffer_reg[0][5]  ( .D(\row2_buffer[1][5] ), .CK(clk), .Q(
        \row2_buffer[0][5] ) );
  DFFQXL \row1_buffer_reg[2][5]  ( .D(\row1_buffer[3][5] ), .CK(clk), .Q(
        \row1_buffer[2][5] ) );
  DFFQXL \row1_buffer_reg[1][5]  ( .D(\row1_buffer[2][5] ), .CK(clk), .Q(
        \row1_buffer[1][5] ) );
  DFFQXL \row3_buffer_reg[2][3]  ( .D(in_pixel[3]), .CK(clk), .Q(
        \row3_buffer[2][3] ) );
  DFFQXL \row3_buffer_reg[1][3]  ( .D(\row3_buffer[2][3] ), .CK(clk), .Q(
        \row3_buffer[1][3] ) );
  DFFQXL \row3_buffer_reg[0][3]  ( .D(\row3_buffer[1][3] ), .CK(clk), .Q(
        \row3_buffer[0][3] ) );
  DFFQXL \row2_buffer_reg[2][3]  ( .D(\row2_buffer[3][3] ), .CK(clk), .Q(
        \row2_buffer[2][3] ) );
  DFFQXL \row2_buffer_reg[1][3]  ( .D(\row2_buffer[2][3] ), .CK(clk), .Q(
        \row2_buffer[1][3] ) );
  DFFQXL \row2_buffer_reg[0][3]  ( .D(\row2_buffer[1][3] ), .CK(clk), .Q(
        \row2_buffer[0][3] ) );
  DFFQXL \row1_buffer_reg[2][3]  ( .D(\row1_buffer[3][3] ), .CK(clk), .Q(
        \row1_buffer[2][3] ) );
  DFFQXL \row1_buffer_reg[1][3]  ( .D(\row1_buffer[2][3] ), .CK(clk), .Q(
        \row1_buffer[1][3] ) );
  DFFQX4 \pixel_00_reg[5]  ( .D(\row1_buffer[0][5] ), .CK(clk), .Q(pixel_00[5]) );
  DFFQX4 \pixel_02_reg[5]  ( .D(\row1_buffer[2][5] ), .CK(clk), .Q(pixel_02[5]) );
  DFFQX4 \pixel_11_reg[5]  ( .D(\row2_buffer[1][5] ), .CK(clk), .Q(pixel_11[5]) );
  DFFQX4 \pixel_20_reg[5]  ( .D(\row3_buffer[0][5] ), .CK(clk), .Q(pixel_20[5]) );
  DFFQX4 \pixel_01_reg[5]  ( .D(\row1_buffer[1][5] ), .CK(clk), .Q(pixel_01[5]) );
  DFFQX4 \pixel_10_reg[5]  ( .D(\row2_buffer[0][5] ), .CK(clk), .Q(pixel_10[5]) );
  DFFQX4 \pixel_12_reg[5]  ( .D(\row2_buffer[2][5] ), .CK(clk), .Q(pixel_12[5]) );
  DFFQX4 \pixel_21_reg[5]  ( .D(\row3_buffer[1][5] ), .CK(clk), .Q(pixel_21[5]) );
  DFFQX4 \pixel_00_reg[3]  ( .D(\row1_buffer[0][3] ), .CK(clk), .Q(pixel_00[3]) );
  DFFQX4 \pixel_02_reg[3]  ( .D(\row1_buffer[2][3] ), .CK(clk), .Q(pixel_02[3]) );
  DFFQX4 \pixel_11_reg[3]  ( .D(\row2_buffer[1][3] ), .CK(clk), .Q(pixel_11[3]) );
  DFFQX4 \pixel_20_reg[3]  ( .D(\row3_buffer[0][3] ), .CK(clk), .Q(pixel_20[3]) );
  DFFQX4 \pixel_01_reg[3]  ( .D(\row1_buffer[1][3] ), .CK(clk), .Q(pixel_01[3]) );
  DFFQX4 \pixel_10_reg[3]  ( .D(\row2_buffer[0][3] ), .CK(clk), .Q(pixel_10[3]) );
  DFFQX4 \pixel_12_reg[3]  ( .D(\row2_buffer[2][3] ), .CK(clk), .Q(pixel_12[3]) );
  DFFQX4 \pixel_21_reg[3]  ( .D(\row3_buffer[1][3] ), .CK(clk), .Q(pixel_21[3]) );
  DFFQX4 \pixel_22_reg[3]  ( .D(\row3_buffer[2][3] ), .CK(clk), .Q(pixel_22[3]) );
  DFFQX4 \pixel_22_reg[5]  ( .D(\row3_buffer[2][5] ), .CK(clk), .Q(pixel_22[5]) );
endmodule


module PE_0_DW_mult_uns_8 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_7 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_6 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_5 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_4 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_3 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0_DW_mult_uns_1 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_0 ( pixel_00, pixel_01, pixel_02, pixel_10, pixel_11, pixel_12, 
        pixel_20, pixel_21, pixel_22, weight_00, weight_01, weight_02, 
        weight_10, weight_11, weight_12, weight_20, weight_21, weight_22, 
        out_pixel_00, out_pixel_01, out_pixel_02, out_pixel_10, out_pixel_11, 
        out_pixel_12, out_pixel_20, out_pixel_21, out_pixel_22, total, clk );
  input [7:0] pixel_00;
  input [7:0] pixel_01;
  input [7:0] pixel_02;
  input [7:0] pixel_10;
  input [7:0] pixel_11;
  input [7:0] pixel_12;
  input [7:0] pixel_20;
  input [7:0] pixel_21;
  input [7:0] pixel_22;
  input [15:0] weight_00;
  input [15:0] weight_01;
  input [15:0] weight_02;
  input [15:0] weight_10;
  input [15:0] weight_11;
  input [15:0] weight_12;
  input [15:0] weight_20;
  input [15:0] weight_21;
  input [15:0] weight_22;
  output [31:0] out_pixel_00;
  output [31:0] out_pixel_01;
  output [31:0] out_pixel_02;
  output [31:0] out_pixel_10;
  output [31:0] out_pixel_11;
  output [31:0] out_pixel_12;
  output [31:0] out_pixel_20;
  output [31:0] out_pixel_21;
  output [31:0] out_pixel_22;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, n1, n2, n3, n4, n5, n6, n7, n8,
         n9;
  assign out_pixel_00[31] = 1'b0;
  assign out_pixel_00[30] = 1'b0;
  assign out_pixel_00[29] = 1'b0;
  assign out_pixel_00[28] = 1'b0;
  assign out_pixel_00[27] = 1'b0;
  assign out_pixel_00[26] = 1'b0;
  assign out_pixel_00[25] = 1'b0;
  assign out_pixel_00[24] = 1'b0;
  assign out_pixel_01[31] = 1'b0;
  assign out_pixel_01[30] = 1'b0;
  assign out_pixel_01[29] = 1'b0;
  assign out_pixel_01[28] = 1'b0;
  assign out_pixel_01[27] = 1'b0;
  assign out_pixel_01[26] = 1'b0;
  assign out_pixel_01[25] = 1'b0;
  assign out_pixel_01[24] = 1'b0;
  assign out_pixel_02[31] = 1'b0;
  assign out_pixel_02[30] = 1'b0;
  assign out_pixel_02[29] = 1'b0;
  assign out_pixel_02[28] = 1'b0;
  assign out_pixel_02[27] = 1'b0;
  assign out_pixel_02[26] = 1'b0;
  assign out_pixel_02[25] = 1'b0;
  assign out_pixel_02[24] = 1'b0;
  assign out_pixel_10[31] = 1'b0;
  assign out_pixel_10[30] = 1'b0;
  assign out_pixel_10[29] = 1'b0;
  assign out_pixel_10[28] = 1'b0;
  assign out_pixel_10[27] = 1'b0;
  assign out_pixel_10[26] = 1'b0;
  assign out_pixel_10[25] = 1'b0;
  assign out_pixel_10[24] = 1'b0;
  assign out_pixel_11[31] = 1'b0;
  assign out_pixel_11[30] = 1'b0;
  assign out_pixel_11[29] = 1'b0;
  assign out_pixel_11[28] = 1'b0;
  assign out_pixel_11[27] = 1'b0;
  assign out_pixel_11[26] = 1'b0;
  assign out_pixel_11[25] = 1'b0;
  assign out_pixel_11[24] = 1'b0;
  assign out_pixel_12[31] = 1'b0;
  assign out_pixel_12[30] = 1'b0;
  assign out_pixel_12[29] = 1'b0;
  assign out_pixel_12[28] = 1'b0;
  assign out_pixel_12[27] = 1'b0;
  assign out_pixel_12[26] = 1'b0;
  assign out_pixel_12[25] = 1'b0;
  assign out_pixel_12[24] = 1'b0;
  assign out_pixel_20[31] = 1'b0;
  assign out_pixel_20[30] = 1'b0;
  assign out_pixel_20[29] = 1'b0;
  assign out_pixel_20[28] = 1'b0;
  assign out_pixel_20[27] = 1'b0;
  assign out_pixel_20[26] = 1'b0;
  assign out_pixel_20[25] = 1'b0;
  assign out_pixel_20[24] = 1'b0;
  assign out_pixel_21[31] = 1'b0;
  assign out_pixel_21[30] = 1'b0;
  assign out_pixel_21[29] = 1'b0;
  assign out_pixel_21[28] = 1'b0;
  assign out_pixel_21[27] = 1'b0;
  assign out_pixel_21[26] = 1'b0;
  assign out_pixel_21[25] = 1'b0;
  assign out_pixel_21[24] = 1'b0;
  assign out_pixel_22[31] = 1'b0;
  assign out_pixel_22[30] = 1'b0;
  assign out_pixel_22[29] = 1'b0;
  assign out_pixel_22[28] = 1'b0;
  assign out_pixel_22[27] = 1'b0;
  assign out_pixel_22[26] = 1'b0;
  assign out_pixel_22[25] = 1'b0;
  assign out_pixel_22[24] = 1'b0;

  PE_0_DW_mult_uns_8 mult_45 ( .a({n1, pixel_22[6:0]}), .b(weight_22), 
        .product({N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192}) );
  PE_0_DW_mult_uns_7 mult_44 ( .a({n2, pixel_21[6:0]}), .b(weight_21), 
        .product({N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, 
        N169, N168}) );
  PE_0_DW_mult_uns_6 mult_43 ( .a({n3, pixel_20[6:0]}), .b(weight_20), 
        .product({N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144}) );
  PE_0_DW_mult_uns_5 mult_42 ( .a({n4, pixel_12[6:0]}), .b(weight_12), 
        .product({N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}) );
  PE_0_DW_mult_uns_4 mult_41 ( .a({n5, pixel_11[6:0]}), .b(weight_11), 
        .product({N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96}) );
  PE_0_DW_mult_uns_3 mult_40 ( .a({n6, pixel_10[6:0]}), .b(weight_10), 
        .product({N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}) );
  PE_0_DW_mult_uns_2 mult_39 ( .a({n7, pixel_02[6:0]}), .b(weight_02), 
        .product({N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48}) );
  PE_0_DW_mult_uns_0 mult_38 ( .a({n8, pixel_01[6:0]}), .b(weight_01), 
        .product({N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24}) );
  PE_0_DW_mult_uns_1 mult_37 ( .a({n9, pixel_00[6:0]}), .b(weight_00), 
        .product({N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  DFFQXL \out_pixel_00_reg[23]  ( .D(N23), .CK(clk), .Q(out_pixel_00[23]) );
  DFFQXL \out_pixel_00_reg[22]  ( .D(N22), .CK(clk), .Q(out_pixel_00[22]) );
  DFFQXL \out_pixel_00_reg[21]  ( .D(N21), .CK(clk), .Q(out_pixel_00[21]) );
  DFFQXL \out_pixel_00_reg[20]  ( .D(N20), .CK(clk), .Q(out_pixel_00[20]) );
  DFFQXL \out_pixel_02_reg[23]  ( .D(N71), .CK(clk), .Q(out_pixel_02[23]) );
  DFFQXL \out_pixel_02_reg[22]  ( .D(N70), .CK(clk), .Q(out_pixel_02[22]) );
  DFFQXL \out_pixel_02_reg[21]  ( .D(N69), .CK(clk), .Q(out_pixel_02[21]) );
  DFFQXL \out_pixel_02_reg[20]  ( .D(N68), .CK(clk), .Q(out_pixel_02[20]) );
  DFFQXL \out_pixel_11_reg[23]  ( .D(N119), .CK(clk), .Q(out_pixel_11[23]) );
  DFFQXL \out_pixel_11_reg[22]  ( .D(N118), .CK(clk), .Q(out_pixel_11[22]) );
  DFFQXL \out_pixel_11_reg[21]  ( .D(N117), .CK(clk), .Q(out_pixel_11[21]) );
  DFFQXL \out_pixel_11_reg[20]  ( .D(N116), .CK(clk), .Q(out_pixel_11[20]) );
  DFFQXL \out_pixel_20_reg[23]  ( .D(N167), .CK(clk), .Q(out_pixel_20[23]) );
  DFFQXL \out_pixel_20_reg[22]  ( .D(N166), .CK(clk), .Q(out_pixel_20[22]) );
  DFFQXL \out_pixel_20_reg[21]  ( .D(N165), .CK(clk), .Q(out_pixel_20[21]) );
  DFFQXL \out_pixel_20_reg[20]  ( .D(N164), .CK(clk), .Q(out_pixel_20[20]) );
  DFFQXL \out_pixel_01_reg[23]  ( .D(N47), .CK(clk), .Q(out_pixel_01[23]) );
  DFFQXL \out_pixel_01_reg[22]  ( .D(N46), .CK(clk), .Q(out_pixel_01[22]) );
  DFFQXL \out_pixel_01_reg[21]  ( .D(N45), .CK(clk), .Q(out_pixel_01[21]) );
  DFFQXL \out_pixel_01_reg[20]  ( .D(N44), .CK(clk), .Q(out_pixel_01[20]) );
  DFFQXL \out_pixel_10_reg[23]  ( .D(N95), .CK(clk), .Q(out_pixel_10[23]) );
  DFFQXL \out_pixel_10_reg[22]  ( .D(N94), .CK(clk), .Q(out_pixel_10[22]) );
  DFFQXL \out_pixel_10_reg[21]  ( .D(N93), .CK(clk), .Q(out_pixel_10[21]) );
  DFFQXL \out_pixel_10_reg[20]  ( .D(N92), .CK(clk), .Q(out_pixel_10[20]) );
  DFFQXL \out_pixel_12_reg[23]  ( .D(N143), .CK(clk), .Q(out_pixel_12[23]) );
  DFFQXL \out_pixel_12_reg[22]  ( .D(N142), .CK(clk), .Q(out_pixel_12[22]) );
  DFFQXL \out_pixel_12_reg[21]  ( .D(N141), .CK(clk), .Q(out_pixel_12[21]) );
  DFFQXL \out_pixel_12_reg[20]  ( .D(N140), .CK(clk), .Q(out_pixel_12[20]) );
  DFFQXL \out_pixel_21_reg[23]  ( .D(N191), .CK(clk), .Q(out_pixel_21[23]) );
  DFFQXL \out_pixel_21_reg[22]  ( .D(N190), .CK(clk), .Q(out_pixel_21[22]) );
  DFFQXL \out_pixel_21_reg[21]  ( .D(N189), .CK(clk), .Q(out_pixel_21[21]) );
  DFFQXL \out_pixel_21_reg[20]  ( .D(N188), .CK(clk), .Q(out_pixel_21[20]) );
  DFFQXL \out_pixel_00_reg[19]  ( .D(N19), .CK(clk), .Q(out_pixel_00[19]) );
  DFFQXL \out_pixel_00_reg[18]  ( .D(N18), .CK(clk), .Q(out_pixel_00[18]) );
  DFFQXL \out_pixel_00_reg[17]  ( .D(N17), .CK(clk), .Q(out_pixel_00[17]) );
  DFFQXL \out_pixel_00_reg[16]  ( .D(N16), .CK(clk), .Q(out_pixel_00[16]) );
  DFFQXL \out_pixel_00_reg[15]  ( .D(N15), .CK(clk), .Q(out_pixel_00[15]) );
  DFFQXL \out_pixel_00_reg[14]  ( .D(N14), .CK(clk), .Q(out_pixel_00[14]) );
  DFFQXL \out_pixel_00_reg[13]  ( .D(N13), .CK(clk), .Q(out_pixel_00[13]) );
  DFFQXL \out_pixel_02_reg[19]  ( .D(N67), .CK(clk), .Q(out_pixel_02[19]) );
  DFFQXL \out_pixel_02_reg[18]  ( .D(N66), .CK(clk), .Q(out_pixel_02[18]) );
  DFFQXL \out_pixel_02_reg[17]  ( .D(N65), .CK(clk), .Q(out_pixel_02[17]) );
  DFFQXL \out_pixel_02_reg[16]  ( .D(N64), .CK(clk), .Q(out_pixel_02[16]) );
  DFFQXL \out_pixel_02_reg[15]  ( .D(N63), .CK(clk), .Q(out_pixel_02[15]) );
  DFFQXL \out_pixel_02_reg[14]  ( .D(N62), .CK(clk), .Q(out_pixel_02[14]) );
  DFFQXL \out_pixel_02_reg[13]  ( .D(N61), .CK(clk), .Q(out_pixel_02[13]) );
  DFFQXL \out_pixel_11_reg[19]  ( .D(N115), .CK(clk), .Q(out_pixel_11[19]) );
  DFFQXL \out_pixel_11_reg[18]  ( .D(N114), .CK(clk), .Q(out_pixel_11[18]) );
  DFFQXL \out_pixel_11_reg[17]  ( .D(N113), .CK(clk), .Q(out_pixel_11[17]) );
  DFFQXL \out_pixel_11_reg[16]  ( .D(N112), .CK(clk), .Q(out_pixel_11[16]) );
  DFFQXL \out_pixel_11_reg[15]  ( .D(N111), .CK(clk), .Q(out_pixel_11[15]) );
  DFFQXL \out_pixel_11_reg[14]  ( .D(N110), .CK(clk), .Q(out_pixel_11[14]) );
  DFFQXL \out_pixel_11_reg[13]  ( .D(N109), .CK(clk), .Q(out_pixel_11[13]) );
  DFFQXL \out_pixel_20_reg[19]  ( .D(N163), .CK(clk), .Q(out_pixel_20[19]) );
  DFFQXL \out_pixel_20_reg[18]  ( .D(N162), .CK(clk), .Q(out_pixel_20[18]) );
  DFFQXL \out_pixel_20_reg[17]  ( .D(N161), .CK(clk), .Q(out_pixel_20[17]) );
  DFFQXL \out_pixel_20_reg[16]  ( .D(N160), .CK(clk), .Q(out_pixel_20[16]) );
  DFFQXL \out_pixel_20_reg[15]  ( .D(N159), .CK(clk), .Q(out_pixel_20[15]) );
  DFFQXL \out_pixel_20_reg[14]  ( .D(N158), .CK(clk), .Q(out_pixel_20[14]) );
  DFFQXL \out_pixel_20_reg[13]  ( .D(N157), .CK(clk), .Q(out_pixel_20[13]) );
  DFFQXL \out_pixel_01_reg[19]  ( .D(N43), .CK(clk), .Q(out_pixel_01[19]) );
  DFFQXL \out_pixel_01_reg[18]  ( .D(N42), .CK(clk), .Q(out_pixel_01[18]) );
  DFFQXL \out_pixel_01_reg[17]  ( .D(N41), .CK(clk), .Q(out_pixel_01[17]) );
  DFFQXL \out_pixel_01_reg[16]  ( .D(N40), .CK(clk), .Q(out_pixel_01[16]) );
  DFFQXL \out_pixel_01_reg[15]  ( .D(N39), .CK(clk), .Q(out_pixel_01[15]) );
  DFFQXL \out_pixel_01_reg[14]  ( .D(N38), .CK(clk), .Q(out_pixel_01[14]) );
  DFFQXL \out_pixel_01_reg[13]  ( .D(N37), .CK(clk), .Q(out_pixel_01[13]) );
  DFFQXL \out_pixel_01_reg[12]  ( .D(N36), .CK(clk), .Q(out_pixel_01[12]) );
  DFFQXL \out_pixel_10_reg[19]  ( .D(N91), .CK(clk), .Q(out_pixel_10[19]) );
  DFFQXL \out_pixel_10_reg[18]  ( .D(N90), .CK(clk), .Q(out_pixel_10[18]) );
  DFFQXL \out_pixel_10_reg[17]  ( .D(N89), .CK(clk), .Q(out_pixel_10[17]) );
  DFFQXL \out_pixel_10_reg[16]  ( .D(N88), .CK(clk), .Q(out_pixel_10[16]) );
  DFFQXL \out_pixel_10_reg[15]  ( .D(N87), .CK(clk), .Q(out_pixel_10[15]) );
  DFFQXL \out_pixel_10_reg[14]  ( .D(N86), .CK(clk), .Q(out_pixel_10[14]) );
  DFFQXL \out_pixel_10_reg[13]  ( .D(N85), .CK(clk), .Q(out_pixel_10[13]) );
  DFFQXL \out_pixel_10_reg[12]  ( .D(N84), .CK(clk), .Q(out_pixel_10[12]) );
  DFFQXL \out_pixel_12_reg[19]  ( .D(N139), .CK(clk), .Q(out_pixel_12[19]) );
  DFFQXL \out_pixel_12_reg[18]  ( .D(N138), .CK(clk), .Q(out_pixel_12[18]) );
  DFFQXL \out_pixel_12_reg[17]  ( .D(N137), .CK(clk), .Q(out_pixel_12[17]) );
  DFFQXL \out_pixel_12_reg[16]  ( .D(N136), .CK(clk), .Q(out_pixel_12[16]) );
  DFFQXL \out_pixel_12_reg[15]  ( .D(N135), .CK(clk), .Q(out_pixel_12[15]) );
  DFFQXL \out_pixel_12_reg[14]  ( .D(N134), .CK(clk), .Q(out_pixel_12[14]) );
  DFFQXL \out_pixel_12_reg[13]  ( .D(N133), .CK(clk), .Q(out_pixel_12[13]) );
  DFFQXL \out_pixel_12_reg[12]  ( .D(N132), .CK(clk), .Q(out_pixel_12[12]) );
  DFFQXL \out_pixel_21_reg[19]  ( .D(N187), .CK(clk), .Q(out_pixel_21[19]) );
  DFFQXL \out_pixel_21_reg[18]  ( .D(N186), .CK(clk), .Q(out_pixel_21[18]) );
  DFFQXL \out_pixel_21_reg[17]  ( .D(N185), .CK(clk), .Q(out_pixel_21[17]) );
  DFFQXL \out_pixel_21_reg[16]  ( .D(N184), .CK(clk), .Q(out_pixel_21[16]) );
  DFFQXL \out_pixel_21_reg[15]  ( .D(N183), .CK(clk), .Q(out_pixel_21[15]) );
  DFFQXL \out_pixel_21_reg[14]  ( .D(N182), .CK(clk), .Q(out_pixel_21[14]) );
  DFFQXL \out_pixel_21_reg[13]  ( .D(N181), .CK(clk), .Q(out_pixel_21[13]) );
  DFFQXL \out_pixel_21_reg[12]  ( .D(N180), .CK(clk), .Q(out_pixel_21[12]) );
  DFFQXL \out_pixel_00_reg[12]  ( .D(N12), .CK(clk), .Q(out_pixel_00[12]) );
  DFFQXL \out_pixel_00_reg[11]  ( .D(N11), .CK(clk), .Q(out_pixel_00[11]) );
  DFFQXL \out_pixel_00_reg[10]  ( .D(N10), .CK(clk), .Q(out_pixel_00[10]) );
  DFFQXL \out_pixel_00_reg[9]  ( .D(N9), .CK(clk), .Q(out_pixel_00[9]) );
  DFFQXL \out_pixel_00_reg[8]  ( .D(N8), .CK(clk), .Q(out_pixel_00[8]) );
  DFFQXL \out_pixel_00_reg[7]  ( .D(N7), .CK(clk), .Q(out_pixel_00[7]) );
  DFFQXL \out_pixel_00_reg[6]  ( .D(N6), .CK(clk), .Q(out_pixel_00[6]) );
  DFFQXL \out_pixel_00_reg[5]  ( .D(N5), .CK(clk), .Q(out_pixel_00[5]) );
  DFFQXL \out_pixel_02_reg[12]  ( .D(N60), .CK(clk), .Q(out_pixel_02[12]) );
  DFFQXL \out_pixel_02_reg[11]  ( .D(N59), .CK(clk), .Q(out_pixel_02[11]) );
  DFFQXL \out_pixel_02_reg[10]  ( .D(N58), .CK(clk), .Q(out_pixel_02[10]) );
  DFFQXL \out_pixel_02_reg[9]  ( .D(N57), .CK(clk), .Q(out_pixel_02[9]) );
  DFFQXL \out_pixel_02_reg[8]  ( .D(N56), .CK(clk), .Q(out_pixel_02[8]) );
  DFFQXL \out_pixel_02_reg[7]  ( .D(N55), .CK(clk), .Q(out_pixel_02[7]) );
  DFFQXL \out_pixel_02_reg[6]  ( .D(N54), .CK(clk), .Q(out_pixel_02[6]) );
  DFFQXL \out_pixel_02_reg[5]  ( .D(N53), .CK(clk), .Q(out_pixel_02[5]) );
  DFFQXL \out_pixel_11_reg[12]  ( .D(N108), .CK(clk), .Q(out_pixel_11[12]) );
  DFFQXL \out_pixel_11_reg[11]  ( .D(N107), .CK(clk), .Q(out_pixel_11[11]) );
  DFFQXL \out_pixel_11_reg[10]  ( .D(N106), .CK(clk), .Q(out_pixel_11[10]) );
  DFFQXL \out_pixel_11_reg[9]  ( .D(N105), .CK(clk), .Q(out_pixel_11[9]) );
  DFFQXL \out_pixel_11_reg[8]  ( .D(N104), .CK(clk), .Q(out_pixel_11[8]) );
  DFFQXL \out_pixel_11_reg[7]  ( .D(N103), .CK(clk), .Q(out_pixel_11[7]) );
  DFFQXL \out_pixel_11_reg[6]  ( .D(N102), .CK(clk), .Q(out_pixel_11[6]) );
  DFFQXL \out_pixel_11_reg[5]  ( .D(N101), .CK(clk), .Q(out_pixel_11[5]) );
  DFFQXL \out_pixel_20_reg[12]  ( .D(N156), .CK(clk), .Q(out_pixel_20[12]) );
  DFFQXL \out_pixel_20_reg[11]  ( .D(N155), .CK(clk), .Q(out_pixel_20[11]) );
  DFFQXL \out_pixel_20_reg[10]  ( .D(N154), .CK(clk), .Q(out_pixel_20[10]) );
  DFFQXL \out_pixel_20_reg[9]  ( .D(N153), .CK(clk), .Q(out_pixel_20[9]) );
  DFFQXL \out_pixel_20_reg[8]  ( .D(N152), .CK(clk), .Q(out_pixel_20[8]) );
  DFFQXL \out_pixel_20_reg[7]  ( .D(N151), .CK(clk), .Q(out_pixel_20[7]) );
  DFFQXL \out_pixel_20_reg[6]  ( .D(N150), .CK(clk), .Q(out_pixel_20[6]) );
  DFFQXL \out_pixel_20_reg[5]  ( .D(N149), .CK(clk), .Q(out_pixel_20[5]) );
  DFFQXL \out_pixel_01_reg[11]  ( .D(N35), .CK(clk), .Q(out_pixel_01[11]) );
  DFFQXL \out_pixel_01_reg[10]  ( .D(N34), .CK(clk), .Q(out_pixel_01[10]) );
  DFFQXL \out_pixel_01_reg[9]  ( .D(N33), .CK(clk), .Q(out_pixel_01[9]) );
  DFFQXL \out_pixel_01_reg[8]  ( .D(N32), .CK(clk), .Q(out_pixel_01[8]) );
  DFFQXL \out_pixel_01_reg[7]  ( .D(N31), .CK(clk), .Q(out_pixel_01[7]) );
  DFFQXL \out_pixel_01_reg[6]  ( .D(N30), .CK(clk), .Q(out_pixel_01[6]) );
  DFFQXL \out_pixel_01_reg[5]  ( .D(N29), .CK(clk), .Q(out_pixel_01[5]) );
  DFFQXL \out_pixel_10_reg[11]  ( .D(N83), .CK(clk), .Q(out_pixel_10[11]) );
  DFFQXL \out_pixel_10_reg[10]  ( .D(N82), .CK(clk), .Q(out_pixel_10[10]) );
  DFFQXL \out_pixel_10_reg[9]  ( .D(N81), .CK(clk), .Q(out_pixel_10[9]) );
  DFFQXL \out_pixel_10_reg[8]  ( .D(N80), .CK(clk), .Q(out_pixel_10[8]) );
  DFFQXL \out_pixel_10_reg[7]  ( .D(N79), .CK(clk), .Q(out_pixel_10[7]) );
  DFFQXL \out_pixel_10_reg[6]  ( .D(N78), .CK(clk), .Q(out_pixel_10[6]) );
  DFFQXL \out_pixel_10_reg[5]  ( .D(N77), .CK(clk), .Q(out_pixel_10[5]) );
  DFFQXL \out_pixel_12_reg[11]  ( .D(N131), .CK(clk), .Q(out_pixel_12[11]) );
  DFFQXL \out_pixel_12_reg[10]  ( .D(N130), .CK(clk), .Q(out_pixel_12[10]) );
  DFFQXL \out_pixel_12_reg[9]  ( .D(N129), .CK(clk), .Q(out_pixel_12[9]) );
  DFFQXL \out_pixel_12_reg[8]  ( .D(N128), .CK(clk), .Q(out_pixel_12[8]) );
  DFFQXL \out_pixel_12_reg[7]  ( .D(N127), .CK(clk), .Q(out_pixel_12[7]) );
  DFFQXL \out_pixel_12_reg[6]  ( .D(N126), .CK(clk), .Q(out_pixel_12[6]) );
  DFFQXL \out_pixel_12_reg[5]  ( .D(N125), .CK(clk), .Q(out_pixel_12[5]) );
  DFFQXL \out_pixel_21_reg[11]  ( .D(N179), .CK(clk), .Q(out_pixel_21[11]) );
  DFFQXL \out_pixel_21_reg[10]  ( .D(N178), .CK(clk), .Q(out_pixel_21[10]) );
  DFFQXL \out_pixel_21_reg[9]  ( .D(N177), .CK(clk), .Q(out_pixel_21[9]) );
  DFFQXL \out_pixel_21_reg[8]  ( .D(N176), .CK(clk), .Q(out_pixel_21[8]) );
  DFFQXL \out_pixel_21_reg[7]  ( .D(N175), .CK(clk), .Q(out_pixel_21[7]) );
  DFFQXL \out_pixel_21_reg[6]  ( .D(N174), .CK(clk), .Q(out_pixel_21[6]) );
  DFFQXL \out_pixel_21_reg[5]  ( .D(N173), .CK(clk), .Q(out_pixel_21[5]) );
  DFFQXL \out_pixel_00_reg[4]  ( .D(N4), .CK(clk), .Q(out_pixel_00[4]) );
  DFFQXL \out_pixel_00_reg[3]  ( .D(N3), .CK(clk), .Q(out_pixel_00[3]) );
  DFFQXL \out_pixel_00_reg[2]  ( .D(N2), .CK(clk), .Q(out_pixel_00[2]) );
  DFFQXL \out_pixel_00_reg[1]  ( .D(N1), .CK(clk), .Q(out_pixel_00[1]) );
  DFFQXL \out_pixel_02_reg[4]  ( .D(N52), .CK(clk), .Q(out_pixel_02[4]) );
  DFFQXL \out_pixel_02_reg[3]  ( .D(N51), .CK(clk), .Q(out_pixel_02[3]) );
  DFFQXL \out_pixel_02_reg[2]  ( .D(N50), .CK(clk), .Q(out_pixel_02[2]) );
  DFFQXL \out_pixel_02_reg[1]  ( .D(N49), .CK(clk), .Q(out_pixel_02[1]) );
  DFFQXL \out_pixel_11_reg[4]  ( .D(N100), .CK(clk), .Q(out_pixel_11[4]) );
  DFFQXL \out_pixel_11_reg[3]  ( .D(N99), .CK(clk), .Q(out_pixel_11[3]) );
  DFFQXL \out_pixel_11_reg[2]  ( .D(N98), .CK(clk), .Q(out_pixel_11[2]) );
  DFFQXL \out_pixel_11_reg[1]  ( .D(N97), .CK(clk), .Q(out_pixel_11[1]) );
  DFFQXL \out_pixel_20_reg[4]  ( .D(N148), .CK(clk), .Q(out_pixel_20[4]) );
  DFFQXL \out_pixel_20_reg[3]  ( .D(N147), .CK(clk), .Q(out_pixel_20[3]) );
  DFFQXL \out_pixel_20_reg[2]  ( .D(N146), .CK(clk), .Q(out_pixel_20[2]) );
  DFFQXL \out_pixel_20_reg[1]  ( .D(N145), .CK(clk), .Q(out_pixel_20[1]) );
  DFFQXL \out_pixel_01_reg[4]  ( .D(N28), .CK(clk), .Q(out_pixel_01[4]) );
  DFFQXL \out_pixel_01_reg[3]  ( .D(N27), .CK(clk), .Q(out_pixel_01[3]) );
  DFFQXL \out_pixel_01_reg[2]  ( .D(N26), .CK(clk), .Q(out_pixel_01[2]) );
  DFFQXL \out_pixel_01_reg[1]  ( .D(N25), .CK(clk), .Q(out_pixel_01[1]) );
  DFFQXL \out_pixel_10_reg[4]  ( .D(N76), .CK(clk), .Q(out_pixel_10[4]) );
  DFFQXL \out_pixel_10_reg[3]  ( .D(N75), .CK(clk), .Q(out_pixel_10[3]) );
  DFFQXL \out_pixel_10_reg[2]  ( .D(N74), .CK(clk), .Q(out_pixel_10[2]) );
  DFFQXL \out_pixel_10_reg[1]  ( .D(N73), .CK(clk), .Q(out_pixel_10[1]) );
  DFFQXL \out_pixel_12_reg[4]  ( .D(N124), .CK(clk), .Q(out_pixel_12[4]) );
  DFFQXL \out_pixel_12_reg[3]  ( .D(N123), .CK(clk), .Q(out_pixel_12[3]) );
  DFFQXL \out_pixel_12_reg[2]  ( .D(N122), .CK(clk), .Q(out_pixel_12[2]) );
  DFFQXL \out_pixel_12_reg[1]  ( .D(N121), .CK(clk), .Q(out_pixel_12[1]) );
  DFFQXL \out_pixel_21_reg[4]  ( .D(N172), .CK(clk), .Q(out_pixel_21[4]) );
  DFFQXL \out_pixel_21_reg[3]  ( .D(N171), .CK(clk), .Q(out_pixel_21[3]) );
  DFFQXL \out_pixel_21_reg[2]  ( .D(N170), .CK(clk), .Q(out_pixel_21[2]) );
  DFFQXL \out_pixel_21_reg[1]  ( .D(N169), .CK(clk), .Q(out_pixel_21[1]) );
  DFFQXL \out_pixel_22_reg[23]  ( .D(N215), .CK(clk), .Q(out_pixel_22[23]) );
  DFFQXL \out_pixel_22_reg[3]  ( .D(N195), .CK(clk), .Q(out_pixel_22[3]) );
  DFFQXL \out_pixel_22_reg[1]  ( .D(N193), .CK(clk), .Q(out_pixel_22[1]) );
  DFFQXL \out_pixel_22_reg[22]  ( .D(N214), .CK(clk), .Q(out_pixel_22[22]) );
  DFFQXL \out_pixel_22_reg[21]  ( .D(N213), .CK(clk), .Q(out_pixel_22[21]) );
  DFFQXL \out_pixel_22_reg[6]  ( .D(N198), .CK(clk), .Q(out_pixel_22[6]) );
  DFFQXL \out_pixel_22_reg[5]  ( .D(N197), .CK(clk), .Q(out_pixel_22[5]) );
  DFFQXL \out_pixel_22_reg[4]  ( .D(N196), .CK(clk), .Q(out_pixel_22[4]) );
  DFFQXL \out_pixel_22_reg[2]  ( .D(N194), .CK(clk), .Q(out_pixel_22[2]) );
  DFFQXL \out_pixel_22_reg[0]  ( .D(N192), .CK(clk), .Q(out_pixel_22[0]) );
  DFFQXL \out_pixel_01_reg[0]  ( .D(N24), .CK(clk), .Q(out_pixel_01[0]) );
  DFFQXL \out_pixel_10_reg[0]  ( .D(N72), .CK(clk), .Q(out_pixel_10[0]) );
  DFFQXL \out_pixel_12_reg[0]  ( .D(N120), .CK(clk), .Q(out_pixel_12[0]) );
  DFFQXL \out_pixel_21_reg[0]  ( .D(N168), .CK(clk), .Q(out_pixel_21[0]) );
  DFFQXL \out_pixel_00_reg[0]  ( .D(N0), .CK(clk), .Q(out_pixel_00[0]) );
  DFFQXL \out_pixel_02_reg[0]  ( .D(N48), .CK(clk), .Q(out_pixel_02[0]) );
  DFFQXL \out_pixel_11_reg[0]  ( .D(N96), .CK(clk), .Q(out_pixel_11[0]) );
  DFFQXL \out_pixel_20_reg[0]  ( .D(N144), .CK(clk), .Q(out_pixel_20[0]) );
  DFFQXL \out_pixel_22_reg[20]  ( .D(N212), .CK(clk), .Q(out_pixel_22[20]) );
  DFFQXL \out_pixel_22_reg[19]  ( .D(N211), .CK(clk), .Q(out_pixel_22[19]) );
  DFFQXL \out_pixel_22_reg[18]  ( .D(N210), .CK(clk), .Q(out_pixel_22[18]) );
  DFFQXL \out_pixel_22_reg[17]  ( .D(N209), .CK(clk), .Q(out_pixel_22[17]) );
  DFFQXL \out_pixel_22_reg[16]  ( .D(N208), .CK(clk), .Q(out_pixel_22[16]) );
  DFFQXL \out_pixel_22_reg[15]  ( .D(N207), .CK(clk), .Q(out_pixel_22[15]) );
  DFFQXL \out_pixel_22_reg[14]  ( .D(N206), .CK(clk), .Q(out_pixel_22[14]) );
  DFFQXL \out_pixel_22_reg[13]  ( .D(N205), .CK(clk), .Q(out_pixel_22[13]) );
  DFFQXL \out_pixel_22_reg[12]  ( .D(N204), .CK(clk), .Q(out_pixel_22[12]) );
  DFFQXL \out_pixel_22_reg[11]  ( .D(N203), .CK(clk), .Q(out_pixel_22[11]) );
  DFFQXL \out_pixel_22_reg[10]  ( .D(N202), .CK(clk), .Q(out_pixel_22[10]) );
  DFFQXL \out_pixel_22_reg[9]  ( .D(N201), .CK(clk), .Q(out_pixel_22[9]) );
  DFFQXL \out_pixel_22_reg[8]  ( .D(N200), .CK(clk), .Q(out_pixel_22[8]) );
  DFFQXL \out_pixel_22_reg[7]  ( .D(N199), .CK(clk), .Q(out_pixel_22[7]) );
  BUFX2 U75 ( .A(pixel_22[7]), .Y(n1) );
  BUFX2 U76 ( .A(pixel_21[7]), .Y(n2) );
  BUFX2 U77 ( .A(pixel_20[7]), .Y(n3) );
  BUFX2 U78 ( .A(pixel_12[7]), .Y(n4) );
  BUFX2 U79 ( .A(pixel_11[7]), .Y(n5) );
  BUFX2 U80 ( .A(pixel_10[7]), .Y(n6) );
  BUFX2 U81 ( .A(pixel_02[7]), .Y(n7) );
  BUFX2 U82 ( .A(pixel_01[7]), .Y(n8) );
  BUFX2 U83 ( .A(pixel_00[7]), .Y(n9) );
endmodule


module PE_3_DW_mult_uns_8 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_7 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_6 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_5 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_4 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_3 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3_DW_mult_uns_1 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_3 ( pixel_00, pixel_01, pixel_02, pixel_10, pixel_11, pixel_12, 
        pixel_20, pixel_21, pixel_22, weight_00, weight_01, weight_02, 
        weight_10, weight_11, weight_12, weight_20, weight_21, weight_22, 
        out_pixel_00, out_pixel_01, out_pixel_02, out_pixel_10, out_pixel_11, 
        out_pixel_12, out_pixel_20, out_pixel_21, out_pixel_22, total, clk );
  input [7:0] pixel_00;
  input [7:0] pixel_01;
  input [7:0] pixel_02;
  input [7:0] pixel_10;
  input [7:0] pixel_11;
  input [7:0] pixel_12;
  input [7:0] pixel_20;
  input [7:0] pixel_21;
  input [7:0] pixel_22;
  input [15:0] weight_00;
  input [15:0] weight_01;
  input [15:0] weight_02;
  input [15:0] weight_10;
  input [15:0] weight_11;
  input [15:0] weight_12;
  input [15:0] weight_20;
  input [15:0] weight_21;
  input [15:0] weight_22;
  output [31:0] out_pixel_00;
  output [31:0] out_pixel_01;
  output [31:0] out_pixel_02;
  output [31:0] out_pixel_10;
  output [31:0] out_pixel_11;
  output [31:0] out_pixel_12;
  output [31:0] out_pixel_20;
  output [31:0] out_pixel_21;
  output [31:0] out_pixel_22;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, n1, n2, n3, n4, n5, n6, n7, n8,
         n9;
  assign out_pixel_00[31] = 1'b0;
  assign out_pixel_00[30] = 1'b0;
  assign out_pixel_00[29] = 1'b0;
  assign out_pixel_00[28] = 1'b0;
  assign out_pixel_00[27] = 1'b0;
  assign out_pixel_00[26] = 1'b0;
  assign out_pixel_00[25] = 1'b0;
  assign out_pixel_00[24] = 1'b0;
  assign out_pixel_01[31] = 1'b0;
  assign out_pixel_01[30] = 1'b0;
  assign out_pixel_01[29] = 1'b0;
  assign out_pixel_01[28] = 1'b0;
  assign out_pixel_01[27] = 1'b0;
  assign out_pixel_01[26] = 1'b0;
  assign out_pixel_01[25] = 1'b0;
  assign out_pixel_01[24] = 1'b0;
  assign out_pixel_02[31] = 1'b0;
  assign out_pixel_02[30] = 1'b0;
  assign out_pixel_02[29] = 1'b0;
  assign out_pixel_02[28] = 1'b0;
  assign out_pixel_02[27] = 1'b0;
  assign out_pixel_02[26] = 1'b0;
  assign out_pixel_02[25] = 1'b0;
  assign out_pixel_02[24] = 1'b0;
  assign out_pixel_10[31] = 1'b0;
  assign out_pixel_10[30] = 1'b0;
  assign out_pixel_10[29] = 1'b0;
  assign out_pixel_10[28] = 1'b0;
  assign out_pixel_10[27] = 1'b0;
  assign out_pixel_10[26] = 1'b0;
  assign out_pixel_10[25] = 1'b0;
  assign out_pixel_10[24] = 1'b0;
  assign out_pixel_11[31] = 1'b0;
  assign out_pixel_11[30] = 1'b0;
  assign out_pixel_11[29] = 1'b0;
  assign out_pixel_11[28] = 1'b0;
  assign out_pixel_11[27] = 1'b0;
  assign out_pixel_11[26] = 1'b0;
  assign out_pixel_11[25] = 1'b0;
  assign out_pixel_11[24] = 1'b0;
  assign out_pixel_12[31] = 1'b0;
  assign out_pixel_12[30] = 1'b0;
  assign out_pixel_12[29] = 1'b0;
  assign out_pixel_12[28] = 1'b0;
  assign out_pixel_12[27] = 1'b0;
  assign out_pixel_12[26] = 1'b0;
  assign out_pixel_12[25] = 1'b0;
  assign out_pixel_12[24] = 1'b0;
  assign out_pixel_20[31] = 1'b0;
  assign out_pixel_20[30] = 1'b0;
  assign out_pixel_20[29] = 1'b0;
  assign out_pixel_20[28] = 1'b0;
  assign out_pixel_20[27] = 1'b0;
  assign out_pixel_20[26] = 1'b0;
  assign out_pixel_20[25] = 1'b0;
  assign out_pixel_20[24] = 1'b0;
  assign out_pixel_21[31] = 1'b0;
  assign out_pixel_21[30] = 1'b0;
  assign out_pixel_21[29] = 1'b0;
  assign out_pixel_21[28] = 1'b0;
  assign out_pixel_21[27] = 1'b0;
  assign out_pixel_21[26] = 1'b0;
  assign out_pixel_21[25] = 1'b0;
  assign out_pixel_21[24] = 1'b0;
  assign out_pixel_22[31] = 1'b0;
  assign out_pixel_22[30] = 1'b0;
  assign out_pixel_22[29] = 1'b0;
  assign out_pixel_22[28] = 1'b0;
  assign out_pixel_22[27] = 1'b0;
  assign out_pixel_22[26] = 1'b0;
  assign out_pixel_22[25] = 1'b0;
  assign out_pixel_22[24] = 1'b0;

  PE_3_DW_mult_uns_8 mult_45 ( .a({n1, pixel_22[6:0]}), .b(weight_22), 
        .product({N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192}) );
  PE_3_DW_mult_uns_7 mult_44 ( .a({n2, pixel_21[6:0]}), .b(weight_21), 
        .product({N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, 
        N169, N168}) );
  PE_3_DW_mult_uns_6 mult_43 ( .a({n3, pixel_20[6:0]}), .b(weight_20), 
        .product({N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144}) );
  PE_3_DW_mult_uns_5 mult_42 ( .a({n4, pixel_12[6:0]}), .b(weight_12), 
        .product({N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}) );
  PE_3_DW_mult_uns_4 mult_41 ( .a({n5, pixel_11[6:0]}), .b(weight_11), 
        .product({N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96}) );
  PE_3_DW_mult_uns_3 mult_40 ( .a({n6, pixel_10[6:0]}), .b(weight_10), 
        .product({N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}) );
  PE_3_DW_mult_uns_2 mult_39 ( .a({n7, pixel_02[6:0]}), .b(weight_02), 
        .product({N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48}) );
  PE_3_DW_mult_uns_0 mult_38 ( .a({n8, pixel_01[6:0]}), .b(weight_01), 
        .product({N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24}) );
  PE_3_DW_mult_uns_1 mult_37 ( .a({n9, pixel_00[6:0]}), .b(weight_00), 
        .product({N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  DFFQXL \out_pixel_00_reg[23]  ( .D(N23), .CK(clk), .Q(out_pixel_00[23]) );
  DFFQXL \out_pixel_00_reg[22]  ( .D(N22), .CK(clk), .Q(out_pixel_00[22]) );
  DFFQXL \out_pixel_00_reg[21]  ( .D(N21), .CK(clk), .Q(out_pixel_00[21]) );
  DFFQXL \out_pixel_00_reg[20]  ( .D(N20), .CK(clk), .Q(out_pixel_00[20]) );
  DFFQXL \out_pixel_02_reg[23]  ( .D(N71), .CK(clk), .Q(out_pixel_02[23]) );
  DFFQXL \out_pixel_02_reg[22]  ( .D(N70), .CK(clk), .Q(out_pixel_02[22]) );
  DFFQXL \out_pixel_02_reg[21]  ( .D(N69), .CK(clk), .Q(out_pixel_02[21]) );
  DFFQXL \out_pixel_02_reg[20]  ( .D(N68), .CK(clk), .Q(out_pixel_02[20]) );
  DFFQXL \out_pixel_11_reg[23]  ( .D(N119), .CK(clk), .Q(out_pixel_11[23]) );
  DFFQXL \out_pixel_11_reg[22]  ( .D(N118), .CK(clk), .Q(out_pixel_11[22]) );
  DFFQXL \out_pixel_11_reg[21]  ( .D(N117), .CK(clk), .Q(out_pixel_11[21]) );
  DFFQXL \out_pixel_11_reg[20]  ( .D(N116), .CK(clk), .Q(out_pixel_11[20]) );
  DFFQXL \out_pixel_20_reg[23]  ( .D(N167), .CK(clk), .Q(out_pixel_20[23]) );
  DFFQXL \out_pixel_20_reg[22]  ( .D(N166), .CK(clk), .Q(out_pixel_20[22]) );
  DFFQXL \out_pixel_20_reg[21]  ( .D(N165), .CK(clk), .Q(out_pixel_20[21]) );
  DFFQXL \out_pixel_20_reg[20]  ( .D(N164), .CK(clk), .Q(out_pixel_20[20]) );
  DFFQXL \out_pixel_01_reg[23]  ( .D(N47), .CK(clk), .Q(out_pixel_01[23]) );
  DFFQXL \out_pixel_01_reg[22]  ( .D(N46), .CK(clk), .Q(out_pixel_01[22]) );
  DFFQXL \out_pixel_01_reg[21]  ( .D(N45), .CK(clk), .Q(out_pixel_01[21]) );
  DFFQXL \out_pixel_01_reg[20]  ( .D(N44), .CK(clk), .Q(out_pixel_01[20]) );
  DFFQXL \out_pixel_10_reg[23]  ( .D(N95), .CK(clk), .Q(out_pixel_10[23]) );
  DFFQXL \out_pixel_10_reg[22]  ( .D(N94), .CK(clk), .Q(out_pixel_10[22]) );
  DFFQXL \out_pixel_10_reg[21]  ( .D(N93), .CK(clk), .Q(out_pixel_10[21]) );
  DFFQXL \out_pixel_10_reg[20]  ( .D(N92), .CK(clk), .Q(out_pixel_10[20]) );
  DFFQXL \out_pixel_12_reg[23]  ( .D(N143), .CK(clk), .Q(out_pixel_12[23]) );
  DFFQXL \out_pixel_12_reg[22]  ( .D(N142), .CK(clk), .Q(out_pixel_12[22]) );
  DFFQXL \out_pixel_12_reg[21]  ( .D(N141), .CK(clk), .Q(out_pixel_12[21]) );
  DFFQXL \out_pixel_12_reg[20]  ( .D(N140), .CK(clk), .Q(out_pixel_12[20]) );
  DFFQXL \out_pixel_21_reg[23]  ( .D(N191), .CK(clk), .Q(out_pixel_21[23]) );
  DFFQXL \out_pixel_21_reg[22]  ( .D(N190), .CK(clk), .Q(out_pixel_21[22]) );
  DFFQXL \out_pixel_21_reg[21]  ( .D(N189), .CK(clk), .Q(out_pixel_21[21]) );
  DFFQXL \out_pixel_21_reg[20]  ( .D(N188), .CK(clk), .Q(out_pixel_21[20]) );
  DFFQXL \out_pixel_00_reg[19]  ( .D(N19), .CK(clk), .Q(out_pixel_00[19]) );
  DFFQXL \out_pixel_00_reg[18]  ( .D(N18), .CK(clk), .Q(out_pixel_00[18]) );
  DFFQXL \out_pixel_00_reg[17]  ( .D(N17), .CK(clk), .Q(out_pixel_00[17]) );
  DFFQXL \out_pixel_00_reg[16]  ( .D(N16), .CK(clk), .Q(out_pixel_00[16]) );
  DFFQXL \out_pixel_00_reg[15]  ( .D(N15), .CK(clk), .Q(out_pixel_00[15]) );
  DFFQXL \out_pixel_00_reg[14]  ( .D(N14), .CK(clk), .Q(out_pixel_00[14]) );
  DFFQXL \out_pixel_00_reg[13]  ( .D(N13), .CK(clk), .Q(out_pixel_00[13]) );
  DFFQXL \out_pixel_02_reg[19]  ( .D(N67), .CK(clk), .Q(out_pixel_02[19]) );
  DFFQXL \out_pixel_02_reg[18]  ( .D(N66), .CK(clk), .Q(out_pixel_02[18]) );
  DFFQXL \out_pixel_02_reg[17]  ( .D(N65), .CK(clk), .Q(out_pixel_02[17]) );
  DFFQXL \out_pixel_02_reg[16]  ( .D(N64), .CK(clk), .Q(out_pixel_02[16]) );
  DFFQXL \out_pixel_02_reg[15]  ( .D(N63), .CK(clk), .Q(out_pixel_02[15]) );
  DFFQXL \out_pixel_02_reg[14]  ( .D(N62), .CK(clk), .Q(out_pixel_02[14]) );
  DFFQXL \out_pixel_02_reg[13]  ( .D(N61), .CK(clk), .Q(out_pixel_02[13]) );
  DFFQXL \out_pixel_11_reg[19]  ( .D(N115), .CK(clk), .Q(out_pixel_11[19]) );
  DFFQXL \out_pixel_11_reg[18]  ( .D(N114), .CK(clk), .Q(out_pixel_11[18]) );
  DFFQXL \out_pixel_11_reg[17]  ( .D(N113), .CK(clk), .Q(out_pixel_11[17]) );
  DFFQXL \out_pixel_11_reg[16]  ( .D(N112), .CK(clk), .Q(out_pixel_11[16]) );
  DFFQXL \out_pixel_11_reg[15]  ( .D(N111), .CK(clk), .Q(out_pixel_11[15]) );
  DFFQXL \out_pixel_11_reg[14]  ( .D(N110), .CK(clk), .Q(out_pixel_11[14]) );
  DFFQXL \out_pixel_11_reg[13]  ( .D(N109), .CK(clk), .Q(out_pixel_11[13]) );
  DFFQXL \out_pixel_20_reg[19]  ( .D(N163), .CK(clk), .Q(out_pixel_20[19]) );
  DFFQXL \out_pixel_20_reg[18]  ( .D(N162), .CK(clk), .Q(out_pixel_20[18]) );
  DFFQXL \out_pixel_20_reg[17]  ( .D(N161), .CK(clk), .Q(out_pixel_20[17]) );
  DFFQXL \out_pixel_20_reg[16]  ( .D(N160), .CK(clk), .Q(out_pixel_20[16]) );
  DFFQXL \out_pixel_20_reg[15]  ( .D(N159), .CK(clk), .Q(out_pixel_20[15]) );
  DFFQXL \out_pixel_20_reg[14]  ( .D(N158), .CK(clk), .Q(out_pixel_20[14]) );
  DFFQXL \out_pixel_20_reg[13]  ( .D(N157), .CK(clk), .Q(out_pixel_20[13]) );
  DFFQXL \out_pixel_01_reg[19]  ( .D(N43), .CK(clk), .Q(out_pixel_01[19]) );
  DFFQXL \out_pixel_01_reg[18]  ( .D(N42), .CK(clk), .Q(out_pixel_01[18]) );
  DFFQXL \out_pixel_01_reg[17]  ( .D(N41), .CK(clk), .Q(out_pixel_01[17]) );
  DFFQXL \out_pixel_01_reg[16]  ( .D(N40), .CK(clk), .Q(out_pixel_01[16]) );
  DFFQXL \out_pixel_01_reg[15]  ( .D(N39), .CK(clk), .Q(out_pixel_01[15]) );
  DFFQXL \out_pixel_01_reg[14]  ( .D(N38), .CK(clk), .Q(out_pixel_01[14]) );
  DFFQXL \out_pixel_01_reg[13]  ( .D(N37), .CK(clk), .Q(out_pixel_01[13]) );
  DFFQXL \out_pixel_01_reg[12]  ( .D(N36), .CK(clk), .Q(out_pixel_01[12]) );
  DFFQXL \out_pixel_10_reg[19]  ( .D(N91), .CK(clk), .Q(out_pixel_10[19]) );
  DFFQXL \out_pixel_10_reg[18]  ( .D(N90), .CK(clk), .Q(out_pixel_10[18]) );
  DFFQXL \out_pixel_10_reg[17]  ( .D(N89), .CK(clk), .Q(out_pixel_10[17]) );
  DFFQXL \out_pixel_10_reg[16]  ( .D(N88), .CK(clk), .Q(out_pixel_10[16]) );
  DFFQXL \out_pixel_10_reg[15]  ( .D(N87), .CK(clk), .Q(out_pixel_10[15]) );
  DFFQXL \out_pixel_10_reg[14]  ( .D(N86), .CK(clk), .Q(out_pixel_10[14]) );
  DFFQXL \out_pixel_10_reg[13]  ( .D(N85), .CK(clk), .Q(out_pixel_10[13]) );
  DFFQXL \out_pixel_10_reg[12]  ( .D(N84), .CK(clk), .Q(out_pixel_10[12]) );
  DFFQXL \out_pixel_12_reg[19]  ( .D(N139), .CK(clk), .Q(out_pixel_12[19]) );
  DFFQXL \out_pixel_12_reg[18]  ( .D(N138), .CK(clk), .Q(out_pixel_12[18]) );
  DFFQXL \out_pixel_12_reg[17]  ( .D(N137), .CK(clk), .Q(out_pixel_12[17]) );
  DFFQXL \out_pixel_12_reg[16]  ( .D(N136), .CK(clk), .Q(out_pixel_12[16]) );
  DFFQXL \out_pixel_12_reg[15]  ( .D(N135), .CK(clk), .Q(out_pixel_12[15]) );
  DFFQXL \out_pixel_12_reg[14]  ( .D(N134), .CK(clk), .Q(out_pixel_12[14]) );
  DFFQXL \out_pixel_12_reg[13]  ( .D(N133), .CK(clk), .Q(out_pixel_12[13]) );
  DFFQXL \out_pixel_12_reg[12]  ( .D(N132), .CK(clk), .Q(out_pixel_12[12]) );
  DFFQXL \out_pixel_21_reg[19]  ( .D(N187), .CK(clk), .Q(out_pixel_21[19]) );
  DFFQXL \out_pixel_21_reg[18]  ( .D(N186), .CK(clk), .Q(out_pixel_21[18]) );
  DFFQXL \out_pixel_21_reg[17]  ( .D(N185), .CK(clk), .Q(out_pixel_21[17]) );
  DFFQXL \out_pixel_21_reg[16]  ( .D(N184), .CK(clk), .Q(out_pixel_21[16]) );
  DFFQXL \out_pixel_21_reg[15]  ( .D(N183), .CK(clk), .Q(out_pixel_21[15]) );
  DFFQXL \out_pixel_21_reg[14]  ( .D(N182), .CK(clk), .Q(out_pixel_21[14]) );
  DFFQXL \out_pixel_21_reg[13]  ( .D(N181), .CK(clk), .Q(out_pixel_21[13]) );
  DFFQXL \out_pixel_21_reg[12]  ( .D(N180), .CK(clk), .Q(out_pixel_21[12]) );
  DFFQXL \out_pixel_00_reg[12]  ( .D(N12), .CK(clk), .Q(out_pixel_00[12]) );
  DFFQXL \out_pixel_00_reg[11]  ( .D(N11), .CK(clk), .Q(out_pixel_00[11]) );
  DFFQXL \out_pixel_00_reg[10]  ( .D(N10), .CK(clk), .Q(out_pixel_00[10]) );
  DFFQXL \out_pixel_00_reg[9]  ( .D(N9), .CK(clk), .Q(out_pixel_00[9]) );
  DFFQXL \out_pixel_00_reg[8]  ( .D(N8), .CK(clk), .Q(out_pixel_00[8]) );
  DFFQXL \out_pixel_00_reg[7]  ( .D(N7), .CK(clk), .Q(out_pixel_00[7]) );
  DFFQXL \out_pixel_00_reg[6]  ( .D(N6), .CK(clk), .Q(out_pixel_00[6]) );
  DFFQXL \out_pixel_00_reg[5]  ( .D(N5), .CK(clk), .Q(out_pixel_00[5]) );
  DFFQXL \out_pixel_02_reg[12]  ( .D(N60), .CK(clk), .Q(out_pixel_02[12]) );
  DFFQXL \out_pixel_02_reg[11]  ( .D(N59), .CK(clk), .Q(out_pixel_02[11]) );
  DFFQXL \out_pixel_02_reg[10]  ( .D(N58), .CK(clk), .Q(out_pixel_02[10]) );
  DFFQXL \out_pixel_02_reg[9]  ( .D(N57), .CK(clk), .Q(out_pixel_02[9]) );
  DFFQXL \out_pixel_02_reg[8]  ( .D(N56), .CK(clk), .Q(out_pixel_02[8]) );
  DFFQXL \out_pixel_02_reg[7]  ( .D(N55), .CK(clk), .Q(out_pixel_02[7]) );
  DFFQXL \out_pixel_02_reg[6]  ( .D(N54), .CK(clk), .Q(out_pixel_02[6]) );
  DFFQXL \out_pixel_02_reg[5]  ( .D(N53), .CK(clk), .Q(out_pixel_02[5]) );
  DFFQXL \out_pixel_11_reg[12]  ( .D(N108), .CK(clk), .Q(out_pixel_11[12]) );
  DFFQXL \out_pixel_11_reg[11]  ( .D(N107), .CK(clk), .Q(out_pixel_11[11]) );
  DFFQXL \out_pixel_11_reg[10]  ( .D(N106), .CK(clk), .Q(out_pixel_11[10]) );
  DFFQXL \out_pixel_11_reg[9]  ( .D(N105), .CK(clk), .Q(out_pixel_11[9]) );
  DFFQXL \out_pixel_11_reg[8]  ( .D(N104), .CK(clk), .Q(out_pixel_11[8]) );
  DFFQXL \out_pixel_11_reg[7]  ( .D(N103), .CK(clk), .Q(out_pixel_11[7]) );
  DFFQXL \out_pixel_11_reg[6]  ( .D(N102), .CK(clk), .Q(out_pixel_11[6]) );
  DFFQXL \out_pixel_11_reg[5]  ( .D(N101), .CK(clk), .Q(out_pixel_11[5]) );
  DFFQXL \out_pixel_20_reg[12]  ( .D(N156), .CK(clk), .Q(out_pixel_20[12]) );
  DFFQXL \out_pixel_20_reg[11]  ( .D(N155), .CK(clk), .Q(out_pixel_20[11]) );
  DFFQXL \out_pixel_20_reg[10]  ( .D(N154), .CK(clk), .Q(out_pixel_20[10]) );
  DFFQXL \out_pixel_20_reg[9]  ( .D(N153), .CK(clk), .Q(out_pixel_20[9]) );
  DFFQXL \out_pixel_20_reg[8]  ( .D(N152), .CK(clk), .Q(out_pixel_20[8]) );
  DFFQXL \out_pixel_20_reg[7]  ( .D(N151), .CK(clk), .Q(out_pixel_20[7]) );
  DFFQXL \out_pixel_20_reg[6]  ( .D(N150), .CK(clk), .Q(out_pixel_20[6]) );
  DFFQXL \out_pixel_20_reg[5]  ( .D(N149), .CK(clk), .Q(out_pixel_20[5]) );
  DFFQXL \out_pixel_01_reg[11]  ( .D(N35), .CK(clk), .Q(out_pixel_01[11]) );
  DFFQXL \out_pixel_01_reg[10]  ( .D(N34), .CK(clk), .Q(out_pixel_01[10]) );
  DFFQXL \out_pixel_01_reg[9]  ( .D(N33), .CK(clk), .Q(out_pixel_01[9]) );
  DFFQXL \out_pixel_01_reg[8]  ( .D(N32), .CK(clk), .Q(out_pixel_01[8]) );
  DFFQXL \out_pixel_01_reg[7]  ( .D(N31), .CK(clk), .Q(out_pixel_01[7]) );
  DFFQXL \out_pixel_01_reg[6]  ( .D(N30), .CK(clk), .Q(out_pixel_01[6]) );
  DFFQXL \out_pixel_01_reg[5]  ( .D(N29), .CK(clk), .Q(out_pixel_01[5]) );
  DFFQXL \out_pixel_10_reg[11]  ( .D(N83), .CK(clk), .Q(out_pixel_10[11]) );
  DFFQXL \out_pixel_10_reg[10]  ( .D(N82), .CK(clk), .Q(out_pixel_10[10]) );
  DFFQXL \out_pixel_10_reg[9]  ( .D(N81), .CK(clk), .Q(out_pixel_10[9]) );
  DFFQXL \out_pixel_10_reg[8]  ( .D(N80), .CK(clk), .Q(out_pixel_10[8]) );
  DFFQXL \out_pixel_10_reg[7]  ( .D(N79), .CK(clk), .Q(out_pixel_10[7]) );
  DFFQXL \out_pixel_10_reg[6]  ( .D(N78), .CK(clk), .Q(out_pixel_10[6]) );
  DFFQXL \out_pixel_10_reg[5]  ( .D(N77), .CK(clk), .Q(out_pixel_10[5]) );
  DFFQXL \out_pixel_12_reg[11]  ( .D(N131), .CK(clk), .Q(out_pixel_12[11]) );
  DFFQXL \out_pixel_12_reg[10]  ( .D(N130), .CK(clk), .Q(out_pixel_12[10]) );
  DFFQXL \out_pixel_12_reg[9]  ( .D(N129), .CK(clk), .Q(out_pixel_12[9]) );
  DFFQXL \out_pixel_12_reg[8]  ( .D(N128), .CK(clk), .Q(out_pixel_12[8]) );
  DFFQXL \out_pixel_12_reg[7]  ( .D(N127), .CK(clk), .Q(out_pixel_12[7]) );
  DFFQXL \out_pixel_12_reg[6]  ( .D(N126), .CK(clk), .Q(out_pixel_12[6]) );
  DFFQXL \out_pixel_12_reg[5]  ( .D(N125), .CK(clk), .Q(out_pixel_12[5]) );
  DFFQXL \out_pixel_21_reg[11]  ( .D(N179), .CK(clk), .Q(out_pixel_21[11]) );
  DFFQXL \out_pixel_21_reg[10]  ( .D(N178), .CK(clk), .Q(out_pixel_21[10]) );
  DFFQXL \out_pixel_21_reg[9]  ( .D(N177), .CK(clk), .Q(out_pixel_21[9]) );
  DFFQXL \out_pixel_21_reg[8]  ( .D(N176), .CK(clk), .Q(out_pixel_21[8]) );
  DFFQXL \out_pixel_21_reg[7]  ( .D(N175), .CK(clk), .Q(out_pixel_21[7]) );
  DFFQXL \out_pixel_21_reg[6]  ( .D(N174), .CK(clk), .Q(out_pixel_21[6]) );
  DFFQXL \out_pixel_21_reg[5]  ( .D(N173), .CK(clk), .Q(out_pixel_21[5]) );
  DFFQXL \out_pixel_00_reg[4]  ( .D(N4), .CK(clk), .Q(out_pixel_00[4]) );
  DFFQXL \out_pixel_00_reg[3]  ( .D(N3), .CK(clk), .Q(out_pixel_00[3]) );
  DFFQXL \out_pixel_00_reg[2]  ( .D(N2), .CK(clk), .Q(out_pixel_00[2]) );
  DFFQXL \out_pixel_00_reg[1]  ( .D(N1), .CK(clk), .Q(out_pixel_00[1]) );
  DFFQXL \out_pixel_02_reg[4]  ( .D(N52), .CK(clk), .Q(out_pixel_02[4]) );
  DFFQXL \out_pixel_02_reg[3]  ( .D(N51), .CK(clk), .Q(out_pixel_02[3]) );
  DFFQXL \out_pixel_02_reg[2]  ( .D(N50), .CK(clk), .Q(out_pixel_02[2]) );
  DFFQXL \out_pixel_02_reg[1]  ( .D(N49), .CK(clk), .Q(out_pixel_02[1]) );
  DFFQXL \out_pixel_11_reg[4]  ( .D(N100), .CK(clk), .Q(out_pixel_11[4]) );
  DFFQXL \out_pixel_11_reg[3]  ( .D(N99), .CK(clk), .Q(out_pixel_11[3]) );
  DFFQXL \out_pixel_11_reg[2]  ( .D(N98), .CK(clk), .Q(out_pixel_11[2]) );
  DFFQXL \out_pixel_11_reg[1]  ( .D(N97), .CK(clk), .Q(out_pixel_11[1]) );
  DFFQXL \out_pixel_20_reg[4]  ( .D(N148), .CK(clk), .Q(out_pixel_20[4]) );
  DFFQXL \out_pixel_20_reg[3]  ( .D(N147), .CK(clk), .Q(out_pixel_20[3]) );
  DFFQXL \out_pixel_20_reg[2]  ( .D(N146), .CK(clk), .Q(out_pixel_20[2]) );
  DFFQXL \out_pixel_20_reg[1]  ( .D(N145), .CK(clk), .Q(out_pixel_20[1]) );
  DFFQXL \out_pixel_01_reg[4]  ( .D(N28), .CK(clk), .Q(out_pixel_01[4]) );
  DFFQXL \out_pixel_01_reg[3]  ( .D(N27), .CK(clk), .Q(out_pixel_01[3]) );
  DFFQXL \out_pixel_01_reg[2]  ( .D(N26), .CK(clk), .Q(out_pixel_01[2]) );
  DFFQXL \out_pixel_01_reg[1]  ( .D(N25), .CK(clk), .Q(out_pixel_01[1]) );
  DFFQXL \out_pixel_10_reg[4]  ( .D(N76), .CK(clk), .Q(out_pixel_10[4]) );
  DFFQXL \out_pixel_10_reg[3]  ( .D(N75), .CK(clk), .Q(out_pixel_10[3]) );
  DFFQXL \out_pixel_10_reg[2]  ( .D(N74), .CK(clk), .Q(out_pixel_10[2]) );
  DFFQXL \out_pixel_10_reg[1]  ( .D(N73), .CK(clk), .Q(out_pixel_10[1]) );
  DFFQXL \out_pixel_12_reg[4]  ( .D(N124), .CK(clk), .Q(out_pixel_12[4]) );
  DFFQXL \out_pixel_12_reg[3]  ( .D(N123), .CK(clk), .Q(out_pixel_12[3]) );
  DFFQXL \out_pixel_12_reg[2]  ( .D(N122), .CK(clk), .Q(out_pixel_12[2]) );
  DFFQXL \out_pixel_12_reg[1]  ( .D(N121), .CK(clk), .Q(out_pixel_12[1]) );
  DFFQXL \out_pixel_21_reg[4]  ( .D(N172), .CK(clk), .Q(out_pixel_21[4]) );
  DFFQXL \out_pixel_21_reg[3]  ( .D(N171), .CK(clk), .Q(out_pixel_21[3]) );
  DFFQXL \out_pixel_21_reg[2]  ( .D(N170), .CK(clk), .Q(out_pixel_21[2]) );
  DFFQXL \out_pixel_21_reg[1]  ( .D(N169), .CK(clk), .Q(out_pixel_21[1]) );
  DFFQXL \out_pixel_22_reg[23]  ( .D(N215), .CK(clk), .Q(out_pixel_22[23]) );
  DFFQXL \out_pixel_22_reg[3]  ( .D(N195), .CK(clk), .Q(out_pixel_22[3]) );
  DFFQXL \out_pixel_22_reg[1]  ( .D(N193), .CK(clk), .Q(out_pixel_22[1]) );
  DFFQXL \out_pixel_22_reg[22]  ( .D(N214), .CK(clk), .Q(out_pixel_22[22]) );
  DFFQXL \out_pixel_22_reg[21]  ( .D(N213), .CK(clk), .Q(out_pixel_22[21]) );
  DFFQXL \out_pixel_22_reg[6]  ( .D(N198), .CK(clk), .Q(out_pixel_22[6]) );
  DFFQXL \out_pixel_22_reg[5]  ( .D(N197), .CK(clk), .Q(out_pixel_22[5]) );
  DFFQXL \out_pixel_22_reg[4]  ( .D(N196), .CK(clk), .Q(out_pixel_22[4]) );
  DFFQXL \out_pixel_22_reg[2]  ( .D(N194), .CK(clk), .Q(out_pixel_22[2]) );
  DFFQXL \out_pixel_22_reg[0]  ( .D(N192), .CK(clk), .Q(out_pixel_22[0]) );
  DFFQXL \out_pixel_01_reg[0]  ( .D(N24), .CK(clk), .Q(out_pixel_01[0]) );
  DFFQXL \out_pixel_10_reg[0]  ( .D(N72), .CK(clk), .Q(out_pixel_10[0]) );
  DFFQXL \out_pixel_12_reg[0]  ( .D(N120), .CK(clk), .Q(out_pixel_12[0]) );
  DFFQXL \out_pixel_21_reg[0]  ( .D(N168), .CK(clk), .Q(out_pixel_21[0]) );
  DFFQXL \out_pixel_00_reg[0]  ( .D(N0), .CK(clk), .Q(out_pixel_00[0]) );
  DFFQXL \out_pixel_02_reg[0]  ( .D(N48), .CK(clk), .Q(out_pixel_02[0]) );
  DFFQXL \out_pixel_11_reg[0]  ( .D(N96), .CK(clk), .Q(out_pixel_11[0]) );
  DFFQXL \out_pixel_20_reg[0]  ( .D(N144), .CK(clk), .Q(out_pixel_20[0]) );
  DFFQXL \out_pixel_22_reg[20]  ( .D(N212), .CK(clk), .Q(out_pixel_22[20]) );
  DFFQXL \out_pixel_22_reg[19]  ( .D(N211), .CK(clk), .Q(out_pixel_22[19]) );
  DFFQXL \out_pixel_22_reg[18]  ( .D(N210), .CK(clk), .Q(out_pixel_22[18]) );
  DFFQXL \out_pixel_22_reg[17]  ( .D(N209), .CK(clk), .Q(out_pixel_22[17]) );
  DFFQXL \out_pixel_22_reg[16]  ( .D(N208), .CK(clk), .Q(out_pixel_22[16]) );
  DFFQXL \out_pixel_22_reg[15]  ( .D(N207), .CK(clk), .Q(out_pixel_22[15]) );
  DFFQXL \out_pixel_22_reg[14]  ( .D(N206), .CK(clk), .Q(out_pixel_22[14]) );
  DFFQXL \out_pixel_22_reg[13]  ( .D(N205), .CK(clk), .Q(out_pixel_22[13]) );
  DFFQXL \out_pixel_22_reg[12]  ( .D(N204), .CK(clk), .Q(out_pixel_22[12]) );
  DFFQXL \out_pixel_22_reg[11]  ( .D(N203), .CK(clk), .Q(out_pixel_22[11]) );
  DFFQXL \out_pixel_22_reg[10]  ( .D(N202), .CK(clk), .Q(out_pixel_22[10]) );
  DFFQXL \out_pixel_22_reg[9]  ( .D(N201), .CK(clk), .Q(out_pixel_22[9]) );
  DFFQXL \out_pixel_22_reg[8]  ( .D(N200), .CK(clk), .Q(out_pixel_22[8]) );
  DFFQXL \out_pixel_22_reg[7]  ( .D(N199), .CK(clk), .Q(out_pixel_22[7]) );
  BUFX2 U75 ( .A(pixel_22[7]), .Y(n1) );
  BUFX2 U76 ( .A(pixel_21[7]), .Y(n2) );
  BUFX2 U77 ( .A(pixel_20[7]), .Y(n3) );
  BUFX2 U78 ( .A(pixel_12[7]), .Y(n4) );
  BUFX2 U79 ( .A(pixel_11[7]), .Y(n5) );
  BUFX2 U80 ( .A(pixel_10[7]), .Y(n6) );
  BUFX2 U81 ( .A(pixel_02[7]), .Y(n7) );
  BUFX2 U82 ( .A(pixel_01[7]), .Y(n8) );
  BUFX2 U83 ( .A(pixel_00[7]), .Y(n9) );
endmodule


module PE_2_DW_mult_uns_8 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_7 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_6 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_5 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_4 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_3 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2_DW_mult_uns_1 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_2 ( pixel_00, pixel_01, pixel_02, pixel_10, pixel_11, pixel_12, 
        pixel_20, pixel_21, pixel_22, weight_00, weight_01, weight_02, 
        weight_10, weight_11, weight_12, weight_20, weight_21, weight_22, 
        out_pixel_00, out_pixel_01, out_pixel_02, out_pixel_10, out_pixel_11, 
        out_pixel_12, out_pixel_20, out_pixel_21, out_pixel_22, total, clk );
  input [7:0] pixel_00;
  input [7:0] pixel_01;
  input [7:0] pixel_02;
  input [7:0] pixel_10;
  input [7:0] pixel_11;
  input [7:0] pixel_12;
  input [7:0] pixel_20;
  input [7:0] pixel_21;
  input [7:0] pixel_22;
  input [15:0] weight_00;
  input [15:0] weight_01;
  input [15:0] weight_02;
  input [15:0] weight_10;
  input [15:0] weight_11;
  input [15:0] weight_12;
  input [15:0] weight_20;
  input [15:0] weight_21;
  input [15:0] weight_22;
  output [31:0] out_pixel_00;
  output [31:0] out_pixel_01;
  output [31:0] out_pixel_02;
  output [31:0] out_pixel_10;
  output [31:0] out_pixel_11;
  output [31:0] out_pixel_12;
  output [31:0] out_pixel_20;
  output [31:0] out_pixel_21;
  output [31:0] out_pixel_22;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, n1, n2, n3, n4, n5, n6, n7, n8,
         n9;
  assign out_pixel_00[31] = 1'b0;
  assign out_pixel_00[30] = 1'b0;
  assign out_pixel_00[29] = 1'b0;
  assign out_pixel_00[28] = 1'b0;
  assign out_pixel_00[27] = 1'b0;
  assign out_pixel_00[26] = 1'b0;
  assign out_pixel_00[25] = 1'b0;
  assign out_pixel_00[24] = 1'b0;
  assign out_pixel_01[31] = 1'b0;
  assign out_pixel_01[30] = 1'b0;
  assign out_pixel_01[29] = 1'b0;
  assign out_pixel_01[28] = 1'b0;
  assign out_pixel_01[27] = 1'b0;
  assign out_pixel_01[26] = 1'b0;
  assign out_pixel_01[25] = 1'b0;
  assign out_pixel_01[24] = 1'b0;
  assign out_pixel_02[31] = 1'b0;
  assign out_pixel_02[30] = 1'b0;
  assign out_pixel_02[29] = 1'b0;
  assign out_pixel_02[28] = 1'b0;
  assign out_pixel_02[27] = 1'b0;
  assign out_pixel_02[26] = 1'b0;
  assign out_pixel_02[25] = 1'b0;
  assign out_pixel_02[24] = 1'b0;
  assign out_pixel_10[31] = 1'b0;
  assign out_pixel_10[30] = 1'b0;
  assign out_pixel_10[29] = 1'b0;
  assign out_pixel_10[28] = 1'b0;
  assign out_pixel_10[27] = 1'b0;
  assign out_pixel_10[26] = 1'b0;
  assign out_pixel_10[25] = 1'b0;
  assign out_pixel_10[24] = 1'b0;
  assign out_pixel_11[31] = 1'b0;
  assign out_pixel_11[30] = 1'b0;
  assign out_pixel_11[29] = 1'b0;
  assign out_pixel_11[28] = 1'b0;
  assign out_pixel_11[27] = 1'b0;
  assign out_pixel_11[26] = 1'b0;
  assign out_pixel_11[25] = 1'b0;
  assign out_pixel_11[24] = 1'b0;
  assign out_pixel_12[31] = 1'b0;
  assign out_pixel_12[30] = 1'b0;
  assign out_pixel_12[29] = 1'b0;
  assign out_pixel_12[28] = 1'b0;
  assign out_pixel_12[27] = 1'b0;
  assign out_pixel_12[26] = 1'b0;
  assign out_pixel_12[25] = 1'b0;
  assign out_pixel_12[24] = 1'b0;
  assign out_pixel_20[31] = 1'b0;
  assign out_pixel_20[30] = 1'b0;
  assign out_pixel_20[29] = 1'b0;
  assign out_pixel_20[28] = 1'b0;
  assign out_pixel_20[27] = 1'b0;
  assign out_pixel_20[26] = 1'b0;
  assign out_pixel_20[25] = 1'b0;
  assign out_pixel_20[24] = 1'b0;
  assign out_pixel_21[31] = 1'b0;
  assign out_pixel_21[30] = 1'b0;
  assign out_pixel_21[29] = 1'b0;
  assign out_pixel_21[28] = 1'b0;
  assign out_pixel_21[27] = 1'b0;
  assign out_pixel_21[26] = 1'b0;
  assign out_pixel_21[25] = 1'b0;
  assign out_pixel_21[24] = 1'b0;
  assign out_pixel_22[31] = 1'b0;
  assign out_pixel_22[30] = 1'b0;
  assign out_pixel_22[29] = 1'b0;
  assign out_pixel_22[28] = 1'b0;
  assign out_pixel_22[27] = 1'b0;
  assign out_pixel_22[26] = 1'b0;
  assign out_pixel_22[25] = 1'b0;
  assign out_pixel_22[24] = 1'b0;

  PE_2_DW_mult_uns_8 mult_45 ( .a({n1, pixel_22[6:0]}), .b(weight_22), 
        .product({N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192}) );
  PE_2_DW_mult_uns_7 mult_44 ( .a({n2, pixel_21[6:0]}), .b(weight_21), 
        .product({N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, 
        N169, N168}) );
  PE_2_DW_mult_uns_6 mult_43 ( .a({n3, pixel_20[6:0]}), .b(weight_20), 
        .product({N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144}) );
  PE_2_DW_mult_uns_5 mult_42 ( .a({n4, pixel_12[6:0]}), .b(weight_12), 
        .product({N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}) );
  PE_2_DW_mult_uns_4 mult_41 ( .a({n5, pixel_11[6:0]}), .b(weight_11), 
        .product({N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96}) );
  PE_2_DW_mult_uns_3 mult_40 ( .a({n6, pixel_10[6:0]}), .b(weight_10), 
        .product({N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}) );
  PE_2_DW_mult_uns_2 mult_39 ( .a({n7, pixel_02[6:0]}), .b(weight_02), 
        .product({N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48}) );
  PE_2_DW_mult_uns_0 mult_38 ( .a({n8, pixel_01[6:0]}), .b(weight_01), 
        .product({N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24}) );
  PE_2_DW_mult_uns_1 mult_37 ( .a({n9, pixel_00[6:0]}), .b(weight_00), 
        .product({N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  DFFQXL \out_pixel_00_reg[23]  ( .D(N23), .CK(clk), .Q(out_pixel_00[23]) );
  DFFQXL \out_pixel_00_reg[22]  ( .D(N22), .CK(clk), .Q(out_pixel_00[22]) );
  DFFQXL \out_pixel_00_reg[21]  ( .D(N21), .CK(clk), .Q(out_pixel_00[21]) );
  DFFQXL \out_pixel_00_reg[20]  ( .D(N20), .CK(clk), .Q(out_pixel_00[20]) );
  DFFQXL \out_pixel_02_reg[23]  ( .D(N71), .CK(clk), .Q(out_pixel_02[23]) );
  DFFQXL \out_pixel_02_reg[22]  ( .D(N70), .CK(clk), .Q(out_pixel_02[22]) );
  DFFQXL \out_pixel_02_reg[21]  ( .D(N69), .CK(clk), .Q(out_pixel_02[21]) );
  DFFQXL \out_pixel_02_reg[20]  ( .D(N68), .CK(clk), .Q(out_pixel_02[20]) );
  DFFQXL \out_pixel_11_reg[23]  ( .D(N119), .CK(clk), .Q(out_pixel_11[23]) );
  DFFQXL \out_pixel_11_reg[22]  ( .D(N118), .CK(clk), .Q(out_pixel_11[22]) );
  DFFQXL \out_pixel_11_reg[21]  ( .D(N117), .CK(clk), .Q(out_pixel_11[21]) );
  DFFQXL \out_pixel_11_reg[20]  ( .D(N116), .CK(clk), .Q(out_pixel_11[20]) );
  DFFQXL \out_pixel_20_reg[23]  ( .D(N167), .CK(clk), .Q(out_pixel_20[23]) );
  DFFQXL \out_pixel_20_reg[22]  ( .D(N166), .CK(clk), .Q(out_pixel_20[22]) );
  DFFQXL \out_pixel_20_reg[21]  ( .D(N165), .CK(clk), .Q(out_pixel_20[21]) );
  DFFQXL \out_pixel_20_reg[20]  ( .D(N164), .CK(clk), .Q(out_pixel_20[20]) );
  DFFQXL \out_pixel_01_reg[23]  ( .D(N47), .CK(clk), .Q(out_pixel_01[23]) );
  DFFQXL \out_pixel_01_reg[22]  ( .D(N46), .CK(clk), .Q(out_pixel_01[22]) );
  DFFQXL \out_pixel_01_reg[21]  ( .D(N45), .CK(clk), .Q(out_pixel_01[21]) );
  DFFQXL \out_pixel_01_reg[20]  ( .D(N44), .CK(clk), .Q(out_pixel_01[20]) );
  DFFQXL \out_pixel_10_reg[23]  ( .D(N95), .CK(clk), .Q(out_pixel_10[23]) );
  DFFQXL \out_pixel_10_reg[22]  ( .D(N94), .CK(clk), .Q(out_pixel_10[22]) );
  DFFQXL \out_pixel_10_reg[21]  ( .D(N93), .CK(clk), .Q(out_pixel_10[21]) );
  DFFQXL \out_pixel_10_reg[20]  ( .D(N92), .CK(clk), .Q(out_pixel_10[20]) );
  DFFQXL \out_pixel_12_reg[23]  ( .D(N143), .CK(clk), .Q(out_pixel_12[23]) );
  DFFQXL \out_pixel_12_reg[22]  ( .D(N142), .CK(clk), .Q(out_pixel_12[22]) );
  DFFQXL \out_pixel_12_reg[21]  ( .D(N141), .CK(clk), .Q(out_pixel_12[21]) );
  DFFQXL \out_pixel_12_reg[20]  ( .D(N140), .CK(clk), .Q(out_pixel_12[20]) );
  DFFQXL \out_pixel_21_reg[23]  ( .D(N191), .CK(clk), .Q(out_pixel_21[23]) );
  DFFQXL \out_pixel_21_reg[22]  ( .D(N190), .CK(clk), .Q(out_pixel_21[22]) );
  DFFQXL \out_pixel_21_reg[21]  ( .D(N189), .CK(clk), .Q(out_pixel_21[21]) );
  DFFQXL \out_pixel_21_reg[20]  ( .D(N188), .CK(clk), .Q(out_pixel_21[20]) );
  DFFQXL \out_pixel_00_reg[19]  ( .D(N19), .CK(clk), .Q(out_pixel_00[19]) );
  DFFQXL \out_pixel_00_reg[18]  ( .D(N18), .CK(clk), .Q(out_pixel_00[18]) );
  DFFQXL \out_pixel_00_reg[17]  ( .D(N17), .CK(clk), .Q(out_pixel_00[17]) );
  DFFQXL \out_pixel_00_reg[16]  ( .D(N16), .CK(clk), .Q(out_pixel_00[16]) );
  DFFQXL \out_pixel_00_reg[15]  ( .D(N15), .CK(clk), .Q(out_pixel_00[15]) );
  DFFQXL \out_pixel_00_reg[14]  ( .D(N14), .CK(clk), .Q(out_pixel_00[14]) );
  DFFQXL \out_pixel_00_reg[13]  ( .D(N13), .CK(clk), .Q(out_pixel_00[13]) );
  DFFQXL \out_pixel_02_reg[19]  ( .D(N67), .CK(clk), .Q(out_pixel_02[19]) );
  DFFQXL \out_pixel_02_reg[18]  ( .D(N66), .CK(clk), .Q(out_pixel_02[18]) );
  DFFQXL \out_pixel_02_reg[17]  ( .D(N65), .CK(clk), .Q(out_pixel_02[17]) );
  DFFQXL \out_pixel_02_reg[16]  ( .D(N64), .CK(clk), .Q(out_pixel_02[16]) );
  DFFQXL \out_pixel_02_reg[15]  ( .D(N63), .CK(clk), .Q(out_pixel_02[15]) );
  DFFQXL \out_pixel_02_reg[14]  ( .D(N62), .CK(clk), .Q(out_pixel_02[14]) );
  DFFQXL \out_pixel_02_reg[13]  ( .D(N61), .CK(clk), .Q(out_pixel_02[13]) );
  DFFQXL \out_pixel_11_reg[19]  ( .D(N115), .CK(clk), .Q(out_pixel_11[19]) );
  DFFQXL \out_pixel_11_reg[18]  ( .D(N114), .CK(clk), .Q(out_pixel_11[18]) );
  DFFQXL \out_pixel_11_reg[17]  ( .D(N113), .CK(clk), .Q(out_pixel_11[17]) );
  DFFQXL \out_pixel_11_reg[16]  ( .D(N112), .CK(clk), .Q(out_pixel_11[16]) );
  DFFQXL \out_pixel_11_reg[15]  ( .D(N111), .CK(clk), .Q(out_pixel_11[15]) );
  DFFQXL \out_pixel_11_reg[14]  ( .D(N110), .CK(clk), .Q(out_pixel_11[14]) );
  DFFQXL \out_pixel_11_reg[13]  ( .D(N109), .CK(clk), .Q(out_pixel_11[13]) );
  DFFQXL \out_pixel_20_reg[19]  ( .D(N163), .CK(clk), .Q(out_pixel_20[19]) );
  DFFQXL \out_pixel_20_reg[18]  ( .D(N162), .CK(clk), .Q(out_pixel_20[18]) );
  DFFQXL \out_pixel_20_reg[17]  ( .D(N161), .CK(clk), .Q(out_pixel_20[17]) );
  DFFQXL \out_pixel_20_reg[16]  ( .D(N160), .CK(clk), .Q(out_pixel_20[16]) );
  DFFQXL \out_pixel_20_reg[15]  ( .D(N159), .CK(clk), .Q(out_pixel_20[15]) );
  DFFQXL \out_pixel_20_reg[14]  ( .D(N158), .CK(clk), .Q(out_pixel_20[14]) );
  DFFQXL \out_pixel_20_reg[13]  ( .D(N157), .CK(clk), .Q(out_pixel_20[13]) );
  DFFQXL \out_pixel_01_reg[19]  ( .D(N43), .CK(clk), .Q(out_pixel_01[19]) );
  DFFQXL \out_pixel_01_reg[18]  ( .D(N42), .CK(clk), .Q(out_pixel_01[18]) );
  DFFQXL \out_pixel_01_reg[17]  ( .D(N41), .CK(clk), .Q(out_pixel_01[17]) );
  DFFQXL \out_pixel_01_reg[16]  ( .D(N40), .CK(clk), .Q(out_pixel_01[16]) );
  DFFQXL \out_pixel_01_reg[15]  ( .D(N39), .CK(clk), .Q(out_pixel_01[15]) );
  DFFQXL \out_pixel_01_reg[14]  ( .D(N38), .CK(clk), .Q(out_pixel_01[14]) );
  DFFQXL \out_pixel_01_reg[13]  ( .D(N37), .CK(clk), .Q(out_pixel_01[13]) );
  DFFQXL \out_pixel_01_reg[12]  ( .D(N36), .CK(clk), .Q(out_pixel_01[12]) );
  DFFQXL \out_pixel_10_reg[19]  ( .D(N91), .CK(clk), .Q(out_pixel_10[19]) );
  DFFQXL \out_pixel_10_reg[18]  ( .D(N90), .CK(clk), .Q(out_pixel_10[18]) );
  DFFQXL \out_pixel_10_reg[17]  ( .D(N89), .CK(clk), .Q(out_pixel_10[17]) );
  DFFQXL \out_pixel_10_reg[16]  ( .D(N88), .CK(clk), .Q(out_pixel_10[16]) );
  DFFQXL \out_pixel_10_reg[15]  ( .D(N87), .CK(clk), .Q(out_pixel_10[15]) );
  DFFQXL \out_pixel_10_reg[14]  ( .D(N86), .CK(clk), .Q(out_pixel_10[14]) );
  DFFQXL \out_pixel_10_reg[13]  ( .D(N85), .CK(clk), .Q(out_pixel_10[13]) );
  DFFQXL \out_pixel_10_reg[12]  ( .D(N84), .CK(clk), .Q(out_pixel_10[12]) );
  DFFQXL \out_pixel_12_reg[19]  ( .D(N139), .CK(clk), .Q(out_pixel_12[19]) );
  DFFQXL \out_pixel_12_reg[18]  ( .D(N138), .CK(clk), .Q(out_pixel_12[18]) );
  DFFQXL \out_pixel_12_reg[17]  ( .D(N137), .CK(clk), .Q(out_pixel_12[17]) );
  DFFQXL \out_pixel_12_reg[16]  ( .D(N136), .CK(clk), .Q(out_pixel_12[16]) );
  DFFQXL \out_pixel_12_reg[15]  ( .D(N135), .CK(clk), .Q(out_pixel_12[15]) );
  DFFQXL \out_pixel_12_reg[14]  ( .D(N134), .CK(clk), .Q(out_pixel_12[14]) );
  DFFQXL \out_pixel_12_reg[13]  ( .D(N133), .CK(clk), .Q(out_pixel_12[13]) );
  DFFQXL \out_pixel_12_reg[12]  ( .D(N132), .CK(clk), .Q(out_pixel_12[12]) );
  DFFQXL \out_pixel_21_reg[19]  ( .D(N187), .CK(clk), .Q(out_pixel_21[19]) );
  DFFQXL \out_pixel_21_reg[18]  ( .D(N186), .CK(clk), .Q(out_pixel_21[18]) );
  DFFQXL \out_pixel_21_reg[17]  ( .D(N185), .CK(clk), .Q(out_pixel_21[17]) );
  DFFQXL \out_pixel_21_reg[16]  ( .D(N184), .CK(clk), .Q(out_pixel_21[16]) );
  DFFQXL \out_pixel_21_reg[15]  ( .D(N183), .CK(clk), .Q(out_pixel_21[15]) );
  DFFQXL \out_pixel_21_reg[14]  ( .D(N182), .CK(clk), .Q(out_pixel_21[14]) );
  DFFQXL \out_pixel_21_reg[13]  ( .D(N181), .CK(clk), .Q(out_pixel_21[13]) );
  DFFQXL \out_pixel_21_reg[12]  ( .D(N180), .CK(clk), .Q(out_pixel_21[12]) );
  DFFQXL \out_pixel_00_reg[12]  ( .D(N12), .CK(clk), .Q(out_pixel_00[12]) );
  DFFQXL \out_pixel_00_reg[11]  ( .D(N11), .CK(clk), .Q(out_pixel_00[11]) );
  DFFQXL \out_pixel_00_reg[10]  ( .D(N10), .CK(clk), .Q(out_pixel_00[10]) );
  DFFQXL \out_pixel_00_reg[9]  ( .D(N9), .CK(clk), .Q(out_pixel_00[9]) );
  DFFQXL \out_pixel_00_reg[8]  ( .D(N8), .CK(clk), .Q(out_pixel_00[8]) );
  DFFQXL \out_pixel_00_reg[7]  ( .D(N7), .CK(clk), .Q(out_pixel_00[7]) );
  DFFQXL \out_pixel_00_reg[6]  ( .D(N6), .CK(clk), .Q(out_pixel_00[6]) );
  DFFQXL \out_pixel_00_reg[5]  ( .D(N5), .CK(clk), .Q(out_pixel_00[5]) );
  DFFQXL \out_pixel_02_reg[12]  ( .D(N60), .CK(clk), .Q(out_pixel_02[12]) );
  DFFQXL \out_pixel_02_reg[11]  ( .D(N59), .CK(clk), .Q(out_pixel_02[11]) );
  DFFQXL \out_pixel_02_reg[10]  ( .D(N58), .CK(clk), .Q(out_pixel_02[10]) );
  DFFQXL \out_pixel_02_reg[9]  ( .D(N57), .CK(clk), .Q(out_pixel_02[9]) );
  DFFQXL \out_pixel_02_reg[8]  ( .D(N56), .CK(clk), .Q(out_pixel_02[8]) );
  DFFQXL \out_pixel_02_reg[7]  ( .D(N55), .CK(clk), .Q(out_pixel_02[7]) );
  DFFQXL \out_pixel_02_reg[6]  ( .D(N54), .CK(clk), .Q(out_pixel_02[6]) );
  DFFQXL \out_pixel_02_reg[5]  ( .D(N53), .CK(clk), .Q(out_pixel_02[5]) );
  DFFQXL \out_pixel_11_reg[12]  ( .D(N108), .CK(clk), .Q(out_pixel_11[12]) );
  DFFQXL \out_pixel_11_reg[11]  ( .D(N107), .CK(clk), .Q(out_pixel_11[11]) );
  DFFQXL \out_pixel_11_reg[10]  ( .D(N106), .CK(clk), .Q(out_pixel_11[10]) );
  DFFQXL \out_pixel_11_reg[9]  ( .D(N105), .CK(clk), .Q(out_pixel_11[9]) );
  DFFQXL \out_pixel_11_reg[8]  ( .D(N104), .CK(clk), .Q(out_pixel_11[8]) );
  DFFQXL \out_pixel_11_reg[7]  ( .D(N103), .CK(clk), .Q(out_pixel_11[7]) );
  DFFQXL \out_pixel_11_reg[6]  ( .D(N102), .CK(clk), .Q(out_pixel_11[6]) );
  DFFQXL \out_pixel_11_reg[5]  ( .D(N101), .CK(clk), .Q(out_pixel_11[5]) );
  DFFQXL \out_pixel_20_reg[12]  ( .D(N156), .CK(clk), .Q(out_pixel_20[12]) );
  DFFQXL \out_pixel_20_reg[11]  ( .D(N155), .CK(clk), .Q(out_pixel_20[11]) );
  DFFQXL \out_pixel_20_reg[10]  ( .D(N154), .CK(clk), .Q(out_pixel_20[10]) );
  DFFQXL \out_pixel_20_reg[9]  ( .D(N153), .CK(clk), .Q(out_pixel_20[9]) );
  DFFQXL \out_pixel_20_reg[8]  ( .D(N152), .CK(clk), .Q(out_pixel_20[8]) );
  DFFQXL \out_pixel_20_reg[7]  ( .D(N151), .CK(clk), .Q(out_pixel_20[7]) );
  DFFQXL \out_pixel_20_reg[6]  ( .D(N150), .CK(clk), .Q(out_pixel_20[6]) );
  DFFQXL \out_pixel_20_reg[5]  ( .D(N149), .CK(clk), .Q(out_pixel_20[5]) );
  DFFQXL \out_pixel_01_reg[11]  ( .D(N35), .CK(clk), .Q(out_pixel_01[11]) );
  DFFQXL \out_pixel_01_reg[10]  ( .D(N34), .CK(clk), .Q(out_pixel_01[10]) );
  DFFQXL \out_pixel_01_reg[9]  ( .D(N33), .CK(clk), .Q(out_pixel_01[9]) );
  DFFQXL \out_pixel_01_reg[8]  ( .D(N32), .CK(clk), .Q(out_pixel_01[8]) );
  DFFQXL \out_pixel_01_reg[7]  ( .D(N31), .CK(clk), .Q(out_pixel_01[7]) );
  DFFQXL \out_pixel_01_reg[6]  ( .D(N30), .CK(clk), .Q(out_pixel_01[6]) );
  DFFQXL \out_pixel_01_reg[5]  ( .D(N29), .CK(clk), .Q(out_pixel_01[5]) );
  DFFQXL \out_pixel_10_reg[11]  ( .D(N83), .CK(clk), .Q(out_pixel_10[11]) );
  DFFQXL \out_pixel_10_reg[10]  ( .D(N82), .CK(clk), .Q(out_pixel_10[10]) );
  DFFQXL \out_pixel_10_reg[9]  ( .D(N81), .CK(clk), .Q(out_pixel_10[9]) );
  DFFQXL \out_pixel_10_reg[8]  ( .D(N80), .CK(clk), .Q(out_pixel_10[8]) );
  DFFQXL \out_pixel_10_reg[7]  ( .D(N79), .CK(clk), .Q(out_pixel_10[7]) );
  DFFQXL \out_pixel_10_reg[6]  ( .D(N78), .CK(clk), .Q(out_pixel_10[6]) );
  DFFQXL \out_pixel_10_reg[5]  ( .D(N77), .CK(clk), .Q(out_pixel_10[5]) );
  DFFQXL \out_pixel_12_reg[11]  ( .D(N131), .CK(clk), .Q(out_pixel_12[11]) );
  DFFQXL \out_pixel_12_reg[10]  ( .D(N130), .CK(clk), .Q(out_pixel_12[10]) );
  DFFQXL \out_pixel_12_reg[9]  ( .D(N129), .CK(clk), .Q(out_pixel_12[9]) );
  DFFQXL \out_pixel_12_reg[8]  ( .D(N128), .CK(clk), .Q(out_pixel_12[8]) );
  DFFQXL \out_pixel_12_reg[7]  ( .D(N127), .CK(clk), .Q(out_pixel_12[7]) );
  DFFQXL \out_pixel_12_reg[6]  ( .D(N126), .CK(clk), .Q(out_pixel_12[6]) );
  DFFQXL \out_pixel_12_reg[5]  ( .D(N125), .CK(clk), .Q(out_pixel_12[5]) );
  DFFQXL \out_pixel_21_reg[11]  ( .D(N179), .CK(clk), .Q(out_pixel_21[11]) );
  DFFQXL \out_pixel_21_reg[10]  ( .D(N178), .CK(clk), .Q(out_pixel_21[10]) );
  DFFQXL \out_pixel_21_reg[9]  ( .D(N177), .CK(clk), .Q(out_pixel_21[9]) );
  DFFQXL \out_pixel_21_reg[8]  ( .D(N176), .CK(clk), .Q(out_pixel_21[8]) );
  DFFQXL \out_pixel_21_reg[7]  ( .D(N175), .CK(clk), .Q(out_pixel_21[7]) );
  DFFQXL \out_pixel_21_reg[6]  ( .D(N174), .CK(clk), .Q(out_pixel_21[6]) );
  DFFQXL \out_pixel_21_reg[5]  ( .D(N173), .CK(clk), .Q(out_pixel_21[5]) );
  DFFQXL \out_pixel_00_reg[4]  ( .D(N4), .CK(clk), .Q(out_pixel_00[4]) );
  DFFQXL \out_pixel_00_reg[3]  ( .D(N3), .CK(clk), .Q(out_pixel_00[3]) );
  DFFQXL \out_pixel_00_reg[2]  ( .D(N2), .CK(clk), .Q(out_pixel_00[2]) );
  DFFQXL \out_pixel_00_reg[1]  ( .D(N1), .CK(clk), .Q(out_pixel_00[1]) );
  DFFQXL \out_pixel_02_reg[4]  ( .D(N52), .CK(clk), .Q(out_pixel_02[4]) );
  DFFQXL \out_pixel_02_reg[3]  ( .D(N51), .CK(clk), .Q(out_pixel_02[3]) );
  DFFQXL \out_pixel_02_reg[2]  ( .D(N50), .CK(clk), .Q(out_pixel_02[2]) );
  DFFQXL \out_pixel_02_reg[1]  ( .D(N49), .CK(clk), .Q(out_pixel_02[1]) );
  DFFQXL \out_pixel_11_reg[4]  ( .D(N100), .CK(clk), .Q(out_pixel_11[4]) );
  DFFQXL \out_pixel_11_reg[3]  ( .D(N99), .CK(clk), .Q(out_pixel_11[3]) );
  DFFQXL \out_pixel_11_reg[2]  ( .D(N98), .CK(clk), .Q(out_pixel_11[2]) );
  DFFQXL \out_pixel_11_reg[1]  ( .D(N97), .CK(clk), .Q(out_pixel_11[1]) );
  DFFQXL \out_pixel_20_reg[4]  ( .D(N148), .CK(clk), .Q(out_pixel_20[4]) );
  DFFQXL \out_pixel_20_reg[3]  ( .D(N147), .CK(clk), .Q(out_pixel_20[3]) );
  DFFQXL \out_pixel_20_reg[2]  ( .D(N146), .CK(clk), .Q(out_pixel_20[2]) );
  DFFQXL \out_pixel_20_reg[1]  ( .D(N145), .CK(clk), .Q(out_pixel_20[1]) );
  DFFQXL \out_pixel_01_reg[4]  ( .D(N28), .CK(clk), .Q(out_pixel_01[4]) );
  DFFQXL \out_pixel_01_reg[3]  ( .D(N27), .CK(clk), .Q(out_pixel_01[3]) );
  DFFQXL \out_pixel_01_reg[2]  ( .D(N26), .CK(clk), .Q(out_pixel_01[2]) );
  DFFQXL \out_pixel_01_reg[1]  ( .D(N25), .CK(clk), .Q(out_pixel_01[1]) );
  DFFQXL \out_pixel_10_reg[4]  ( .D(N76), .CK(clk), .Q(out_pixel_10[4]) );
  DFFQXL \out_pixel_10_reg[3]  ( .D(N75), .CK(clk), .Q(out_pixel_10[3]) );
  DFFQXL \out_pixel_10_reg[2]  ( .D(N74), .CK(clk), .Q(out_pixel_10[2]) );
  DFFQXL \out_pixel_10_reg[1]  ( .D(N73), .CK(clk), .Q(out_pixel_10[1]) );
  DFFQXL \out_pixel_12_reg[4]  ( .D(N124), .CK(clk), .Q(out_pixel_12[4]) );
  DFFQXL \out_pixel_12_reg[3]  ( .D(N123), .CK(clk), .Q(out_pixel_12[3]) );
  DFFQXL \out_pixel_12_reg[2]  ( .D(N122), .CK(clk), .Q(out_pixel_12[2]) );
  DFFQXL \out_pixel_12_reg[1]  ( .D(N121), .CK(clk), .Q(out_pixel_12[1]) );
  DFFQXL \out_pixel_21_reg[4]  ( .D(N172), .CK(clk), .Q(out_pixel_21[4]) );
  DFFQXL \out_pixel_21_reg[3]  ( .D(N171), .CK(clk), .Q(out_pixel_21[3]) );
  DFFQXL \out_pixel_21_reg[2]  ( .D(N170), .CK(clk), .Q(out_pixel_21[2]) );
  DFFQXL \out_pixel_21_reg[1]  ( .D(N169), .CK(clk), .Q(out_pixel_21[1]) );
  DFFQXL \out_pixel_22_reg[23]  ( .D(N215), .CK(clk), .Q(out_pixel_22[23]) );
  DFFQXL \out_pixel_22_reg[3]  ( .D(N195), .CK(clk), .Q(out_pixel_22[3]) );
  DFFQXL \out_pixel_22_reg[1]  ( .D(N193), .CK(clk), .Q(out_pixel_22[1]) );
  DFFQXL \out_pixel_22_reg[22]  ( .D(N214), .CK(clk), .Q(out_pixel_22[22]) );
  DFFQXL \out_pixel_22_reg[21]  ( .D(N213), .CK(clk), .Q(out_pixel_22[21]) );
  DFFQXL \out_pixel_22_reg[6]  ( .D(N198), .CK(clk), .Q(out_pixel_22[6]) );
  DFFQXL \out_pixel_22_reg[5]  ( .D(N197), .CK(clk), .Q(out_pixel_22[5]) );
  DFFQXL \out_pixel_22_reg[4]  ( .D(N196), .CK(clk), .Q(out_pixel_22[4]) );
  DFFQXL \out_pixel_22_reg[2]  ( .D(N194), .CK(clk), .Q(out_pixel_22[2]) );
  DFFQXL \out_pixel_22_reg[0]  ( .D(N192), .CK(clk), .Q(out_pixel_22[0]) );
  DFFQXL \out_pixel_01_reg[0]  ( .D(N24), .CK(clk), .Q(out_pixel_01[0]) );
  DFFQXL \out_pixel_10_reg[0]  ( .D(N72), .CK(clk), .Q(out_pixel_10[0]) );
  DFFQXL \out_pixel_12_reg[0]  ( .D(N120), .CK(clk), .Q(out_pixel_12[0]) );
  DFFQXL \out_pixel_21_reg[0]  ( .D(N168), .CK(clk), .Q(out_pixel_21[0]) );
  DFFQXL \out_pixel_00_reg[0]  ( .D(N0), .CK(clk), .Q(out_pixel_00[0]) );
  DFFQXL \out_pixel_02_reg[0]  ( .D(N48), .CK(clk), .Q(out_pixel_02[0]) );
  DFFQXL \out_pixel_11_reg[0]  ( .D(N96), .CK(clk), .Q(out_pixel_11[0]) );
  DFFQXL \out_pixel_20_reg[0]  ( .D(N144), .CK(clk), .Q(out_pixel_20[0]) );
  DFFQXL \out_pixel_22_reg[20]  ( .D(N212), .CK(clk), .Q(out_pixel_22[20]) );
  DFFQXL \out_pixel_22_reg[19]  ( .D(N211), .CK(clk), .Q(out_pixel_22[19]) );
  DFFQXL \out_pixel_22_reg[18]  ( .D(N210), .CK(clk), .Q(out_pixel_22[18]) );
  DFFQXL \out_pixel_22_reg[17]  ( .D(N209), .CK(clk), .Q(out_pixel_22[17]) );
  DFFQXL \out_pixel_22_reg[16]  ( .D(N208), .CK(clk), .Q(out_pixel_22[16]) );
  DFFQXL \out_pixel_22_reg[15]  ( .D(N207), .CK(clk), .Q(out_pixel_22[15]) );
  DFFQXL \out_pixel_22_reg[14]  ( .D(N206), .CK(clk), .Q(out_pixel_22[14]) );
  DFFQXL \out_pixel_22_reg[13]  ( .D(N205), .CK(clk), .Q(out_pixel_22[13]) );
  DFFQXL \out_pixel_22_reg[12]  ( .D(N204), .CK(clk), .Q(out_pixel_22[12]) );
  DFFQXL \out_pixel_22_reg[11]  ( .D(N203), .CK(clk), .Q(out_pixel_22[11]) );
  DFFQXL \out_pixel_22_reg[10]  ( .D(N202), .CK(clk), .Q(out_pixel_22[10]) );
  DFFQXL \out_pixel_22_reg[9]  ( .D(N201), .CK(clk), .Q(out_pixel_22[9]) );
  DFFQXL \out_pixel_22_reg[8]  ( .D(N200), .CK(clk), .Q(out_pixel_22[8]) );
  DFFQXL \out_pixel_22_reg[7]  ( .D(N199), .CK(clk), .Q(out_pixel_22[7]) );
  BUFX2 U75 ( .A(pixel_22[7]), .Y(n1) );
  BUFX2 U76 ( .A(pixel_21[7]), .Y(n2) );
  BUFX2 U77 ( .A(pixel_20[7]), .Y(n3) );
  BUFX2 U78 ( .A(pixel_12[7]), .Y(n4) );
  BUFX2 U79 ( .A(pixel_11[7]), .Y(n5) );
  BUFX2 U80 ( .A(pixel_10[7]), .Y(n6) );
  BUFX2 U81 ( .A(pixel_02[7]), .Y(n7) );
  BUFX2 U82 ( .A(pixel_01[7]), .Y(n8) );
  BUFX2 U83 ( .A(pixel_00[7]), .Y(n9) );
endmodule


module PE_1_DW_mult_uns_8 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_7 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_6 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_5 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_4 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_3 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1_DW_mult_uns_1 ( a, b, product );
  input [7:0] a;
  input [15:0] b;
  output [23:0] product;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n52, n53, n54, n55,
         n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;

  ADDFX1 U27 ( .A(n54), .B(n50), .CI(n27), .CO(n26), .S(product[22]) );
  ADDFX1 U28 ( .A(n57), .B(n55), .CI(n28), .CO(n27), .S(product[21]) );
  ADDFX1 U29 ( .A(n58), .B(n62), .CI(n29), .CO(n28), .S(product[20]) );
  ADDFX1 U30 ( .A(n63), .B(n67), .CI(n30), .CO(n29), .S(product[19]) );
  ADDFX1 U31 ( .A(n68), .B(n74), .CI(n31), .CO(n30), .S(product[18]) );
  ADDFX1 U32 ( .A(n75), .B(n80), .CI(n32), .CO(n31), .S(product[17]) );
  ADDFX1 U33 ( .A(n81), .B(n85), .CI(n33), .CO(n32), .S(product[16]) );
  ADDFX1 U34 ( .A(n86), .B(n90), .CI(n34), .CO(n33), .S(product[15]) );
  ADDFX1 U35 ( .A(n91), .B(n95), .CI(n35), .CO(n34), .S(product[14]) );
  ADDFX1 U36 ( .A(n96), .B(n100), .CI(n36), .CO(n35), .S(product[13]) );
  ADDFX1 U37 ( .A(n101), .B(n105), .CI(n37), .CO(n36), .S(product[12]) );
  ADDFX1 U38 ( .A(n106), .B(n110), .CI(n38), .CO(n37), .S(product[11]) );
  ADDFX1 U39 ( .A(n111), .B(n115), .CI(n39), .CO(n38), .S(product[10]) );
  ADDFX1 U40 ( .A(n116), .B(n120), .CI(n40), .CO(n39), .S(product[9]) );
  ADDFX1 U41 ( .A(n121), .B(n125), .CI(n41), .CO(n40), .S(product[8]) );
  ADDFX1 U42 ( .A(n126), .B(n130), .CI(n42), .CO(n41), .S(product[7]) );
  ADDFX1 U43 ( .A(n131), .B(n132), .CI(n43), .CO(n42), .S(product[6]) );
  ADDFX1 U44 ( .A(n133), .B(n136), .CI(n44), .CO(n43), .S(product[5]) );
  ADDFX1 U45 ( .A(n137), .B(n138), .CI(n45), .CO(n44), .S(product[4]) );
  ADDFX1 U46 ( .A(n139), .B(n142), .CI(n46), .CO(n45), .S(product[3]) );
  ADDFX1 U47 ( .A(n226), .B(n210), .CI(n47), .CO(n46), .S(product[2]) );
  ADDHX1 U48 ( .A(n143), .B(n227), .CO(n47), .S(product[1]) );
  ADDFX1 U50 ( .A(n158), .B(n52), .CI(n53), .CO(n49), .S(n50) );
  CMPR42X1 U52 ( .A(n408), .B(n145), .C(n175), .D(n159), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U53 ( .A(n60), .B(n176), .C(n160), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U55 ( .A(n177), .B(n161), .C(n65), .D(n69), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFX1 U56 ( .A(n146), .B(n407), .CI(n193), .CO(n64), .S(n65) );
  CMPR42X1 U57 ( .A(n178), .B(n162), .C(n70), .D(n76), .ICI(n73), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFX1 U58 ( .A(n78), .B(n147), .CI(n194), .CO(n69), .S(n70) );
  CMPR42X1 U60 ( .A(n179), .B(n163), .C(n77), .D(n82), .ICI(n79), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFX1 U61 ( .A(n411), .B(n78), .CI(n195), .CO(n76), .S(n77) );
  CMPR42X1 U63 ( .A(n180), .B(n164), .C(n87), .D(n83), .ICI(n84), .S(n81), 
        .ICO(n79), .CO(n80) );
  ADDFX1 U64 ( .A(n212), .B(n148), .CI(n196), .CO(n82), .S(n83) );
  CMPR42X1 U65 ( .A(n181), .B(n165), .C(n92), .D(n88), .ICI(n89), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFX1 U66 ( .A(n213), .B(n149), .CI(n197), .CO(n87), .S(n88) );
  CMPR42X1 U67 ( .A(n182), .B(n166), .C(n97), .D(n93), .ICI(n94), .S(n91), 
        .ICO(n89), .CO(n90) );
  ADDFX1 U68 ( .A(n214), .B(n150), .CI(n198), .CO(n92), .S(n93) );
  CMPR42X1 U69 ( .A(n183), .B(n167), .C(n102), .D(n98), .ICI(n99), .S(n96), 
        .ICO(n94), .CO(n95) );
  ADDFX1 U70 ( .A(n215), .B(n151), .CI(n199), .CO(n97), .S(n98) );
  CMPR42X1 U71 ( .A(n184), .B(n168), .C(n107), .D(n103), .ICI(n104), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDFX1 U72 ( .A(n216), .B(n152), .CI(n200), .CO(n102), .S(n103) );
  CMPR42X1 U73 ( .A(n185), .B(n169), .C(n112), .D(n108), .ICI(n109), .S(n106), 
        .ICO(n104), .CO(n105) );
  ADDFX1 U74 ( .A(n217), .B(n153), .CI(n201), .CO(n107), .S(n108) );
  CMPR42X1 U75 ( .A(n186), .B(n170), .C(n117), .D(n113), .ICI(n114), .S(n111), 
        .ICO(n109), .CO(n110) );
  ADDFX1 U76 ( .A(n218), .B(n154), .CI(n202), .CO(n112), .S(n113) );
  CMPR42X1 U77 ( .A(n187), .B(n171), .C(n122), .D(n118), .ICI(n119), .S(n116), 
        .ICO(n114), .CO(n115) );
  ADDFX1 U78 ( .A(n219), .B(n155), .CI(n203), .CO(n117), .S(n118) );
  CMPR42X1 U79 ( .A(n188), .B(n172), .C(n127), .D(n124), .ICI(n123), .S(n121), 
        .ICO(n119), .CO(n120) );
  ADDFX1 U80 ( .A(n220), .B(n156), .CI(n204), .CO(n122), .S(n123) );
  CMPR42X1 U81 ( .A(n205), .B(n173), .C(n189), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDHX1 U82 ( .A(n221), .B(n140), .CO(n127), .S(n128) );
  CMPR42X1 U83 ( .A(n174), .B(n222), .C(n206), .D(n190), .ICI(n134), .S(n131), 
        .ICO(n129), .CO(n130) );
  ADDFX1 U84 ( .A(n191), .B(n207), .CI(n135), .CO(n132), .S(n133) );
  ADDHX1 U85 ( .A(n223), .B(n141), .CO(n134), .S(n135) );
  ADDFX1 U86 ( .A(n224), .B(n192), .CI(n208), .CO(n136), .S(n137) );
  ADDHX1 U87 ( .A(n225), .B(n209), .CO(n138), .S(n139) );
  INVX4 U299 ( .A(a[7]), .Y(n405) );
  INVX4 U300 ( .A(a[7]), .Y(n404) );
  BUFX2 U301 ( .A(a[7]), .Y(n406) );
  INVX5 U302 ( .A(a[3]), .Y(n410) );
  INVX5 U303 ( .A(a[5]), .Y(n409) );
  INVX5 U304 ( .A(a[1]), .Y(n411) );
  INVX4 U305 ( .A(a[0]), .Y(n412) );
  BUFX5 U306 ( .A(n420), .Y(n403) );
  XOR2X1 U307 ( .A(a[6]), .B(n409), .Y(n420) );
  BUFX5 U308 ( .A(n455), .Y(n401) );
  XOR2X1 U309 ( .A(a[4]), .B(n410), .Y(n455) );
  BUFX5 U310 ( .A(n437), .Y(n399) );
  XOR2X1 U311 ( .A(a[2]), .B(n411), .Y(n437) );
  CLKBUFX4 U312 ( .A(n457), .Y(n400) );
  NAND2X2 U313 ( .A(n401), .B(n490), .Y(n457) );
  CLKBUFX4 U314 ( .A(n439), .Y(n398) );
  NAND2X2 U315 ( .A(n399), .B(n489), .Y(n439) );
  CLKBUFX4 U316 ( .A(n419), .Y(n402) );
  NAND2X2 U317 ( .A(n403), .B(n491), .Y(n419) );
  CLKBUFX4 U318 ( .A(n421), .Y(n397) );
  NAND2X2 U319 ( .A(a[1]), .B(n412), .Y(n421) );
  INVX2 U320 ( .A(b[0]), .Y(n413) );
  INVX2 U321 ( .A(n78), .Y(n407) );
  INVX2 U322 ( .A(n60), .Y(n408) );
  XOR2X1 U323 ( .A(n414), .B(n415), .Y(product[23]) );
  XOR2X1 U324 ( .A(n52), .B(n416), .Y(n415) );
  XNOR2X1 U325 ( .A(n49), .B(n26), .Y(n416) );
  XOR2X1 U326 ( .A(n417), .B(n418), .Y(n414) );
  AND2X1 U327 ( .A(b[15]), .B(n406), .Y(n418) );
  OAI2BB1X1 U328 ( .A0N(n402), .A1N(n403), .B0(n406), .Y(n417) );
  NOR2X1 U329 ( .A(n413), .B(n412), .Y(product[0]) );
  CLKNAND2X2 U330 ( .A(b[9]), .B(a[7]), .Y(n78) );
  CLKNAND2X2 U331 ( .A(b[12]), .B(a[7]), .Y(n60) );
  CLKNAND2X2 U332 ( .A(b[14]), .B(a[7]), .Y(n52) );
  OAI22X1 U333 ( .A0(b[0]), .A1(n397), .B0(n422), .B1(n412), .Y(n227) );
  OAI22X1 U334 ( .A0(n422), .A1(n397), .B0(n423), .B1(n412), .Y(n226) );
  XOR2X1 U335 ( .A(b[1]), .B(n411), .Y(n422) );
  OAI22X1 U336 ( .A0(n423), .A1(n397), .B0(n424), .B1(n412), .Y(n225) );
  XOR2X1 U337 ( .A(b[2]), .B(n411), .Y(n423) );
  OAI22X1 U338 ( .A0(n424), .A1(n397), .B0(n425), .B1(n412), .Y(n224) );
  XOR2X1 U339 ( .A(b[3]), .B(n411), .Y(n424) );
  OAI22X1 U340 ( .A0(n425), .A1(n397), .B0(n426), .B1(n412), .Y(n223) );
  XOR2X1 U341 ( .A(b[4]), .B(n411), .Y(n425) );
  OAI22X1 U342 ( .A0(n426), .A1(n397), .B0(n427), .B1(n412), .Y(n222) );
  XOR2X1 U343 ( .A(b[5]), .B(n411), .Y(n426) );
  OAI22X1 U344 ( .A0(n427), .A1(n397), .B0(n428), .B1(n412), .Y(n221) );
  XOR2X1 U345 ( .A(b[6]), .B(n411), .Y(n427) );
  OAI22X1 U346 ( .A0(n428), .A1(n397), .B0(n429), .B1(n412), .Y(n220) );
  XOR2X1 U347 ( .A(b[7]), .B(n411), .Y(n428) );
  OAI22X1 U348 ( .A0(n429), .A1(n397), .B0(n430), .B1(n412), .Y(n219) );
  XOR2X1 U349 ( .A(b[8]), .B(n411), .Y(n429) );
  OAI22X1 U350 ( .A0(n430), .A1(n397), .B0(n431), .B1(n412), .Y(n218) );
  XOR2X1 U351 ( .A(b[9]), .B(n411), .Y(n430) );
  OAI22X1 U352 ( .A0(n431), .A1(n397), .B0(n432), .B1(n412), .Y(n217) );
  XOR2X1 U353 ( .A(b[10]), .B(n411), .Y(n431) );
  OAI22X1 U354 ( .A0(n432), .A1(n397), .B0(n433), .B1(n412), .Y(n216) );
  XOR2X1 U355 ( .A(b[11]), .B(n411), .Y(n432) );
  OAI22X1 U356 ( .A0(n433), .A1(n397), .B0(n434), .B1(n412), .Y(n215) );
  XOR2X1 U357 ( .A(b[12]), .B(n411), .Y(n433) );
  OAI22X1 U358 ( .A0(n434), .A1(n397), .B0(n435), .B1(n412), .Y(n214) );
  XOR2X1 U359 ( .A(b[13]), .B(n411), .Y(n434) );
  OAI22X1 U360 ( .A0(n435), .A1(n397), .B0(n436), .B1(n412), .Y(n213) );
  XOR2X1 U361 ( .A(b[14]), .B(n411), .Y(n435) );
  OAI22X1 U362 ( .A0(n436), .A1(n397), .B0(n412), .B1(n411), .Y(n212) );
  XOR2X1 U363 ( .A(b[15]), .B(n411), .Y(n436) );
  NOR2X1 U364 ( .A(n413), .B(n399), .Y(n210) );
  OAI22X1 U365 ( .A0(n438), .A1(n398), .B0(n399), .B1(n440), .Y(n209) );
  XOR2X1 U366 ( .A(n413), .B(a[3]), .Y(n438) );
  OAI22X1 U367 ( .A0(n440), .A1(n398), .B0(n399), .B1(n441), .Y(n208) );
  XOR2X1 U368 ( .A(b[1]), .B(n410), .Y(n440) );
  OAI22X1 U369 ( .A0(n441), .A1(n398), .B0(n399), .B1(n442), .Y(n207) );
  XOR2X1 U370 ( .A(b[2]), .B(n410), .Y(n441) );
  OAI22X1 U371 ( .A0(n442), .A1(n398), .B0(n399), .B1(n443), .Y(n206) );
  XOR2X1 U372 ( .A(b[3]), .B(n410), .Y(n442) );
  OAI22X1 U373 ( .A0(n443), .A1(n398), .B0(n399), .B1(n444), .Y(n205) );
  XOR2X1 U374 ( .A(b[4]), .B(n410), .Y(n443) );
  OAI22X1 U375 ( .A0(n444), .A1(n398), .B0(n399), .B1(n445), .Y(n204) );
  XOR2X1 U376 ( .A(b[5]), .B(n410), .Y(n444) );
  OAI22X1 U377 ( .A0(n445), .A1(n398), .B0(n399), .B1(n446), .Y(n203) );
  XOR2X1 U378 ( .A(b[6]), .B(n410), .Y(n445) );
  OAI22X1 U379 ( .A0(n446), .A1(n398), .B0(n399), .B1(n447), .Y(n202) );
  XOR2X1 U380 ( .A(b[7]), .B(n410), .Y(n446) );
  OAI22X1 U381 ( .A0(n447), .A1(n398), .B0(n399), .B1(n448), .Y(n201) );
  XOR2X1 U382 ( .A(b[8]), .B(n410), .Y(n447) );
  OAI22X1 U383 ( .A0(n448), .A1(n398), .B0(n399), .B1(n449), .Y(n200) );
  XOR2X1 U384 ( .A(b[9]), .B(n410), .Y(n448) );
  OAI22X1 U385 ( .A0(n449), .A1(n398), .B0(n399), .B1(n450), .Y(n199) );
  XOR2X1 U386 ( .A(b[10]), .B(n410), .Y(n449) );
  OAI22X1 U387 ( .A0(n450), .A1(n398), .B0(n399), .B1(n451), .Y(n198) );
  XOR2X1 U388 ( .A(b[11]), .B(n410), .Y(n450) );
  OAI22X1 U389 ( .A0(n451), .A1(n398), .B0(n399), .B1(n452), .Y(n197) );
  XOR2X1 U390 ( .A(b[12]), .B(n410), .Y(n451) );
  OAI22X1 U391 ( .A0(n452), .A1(n398), .B0(n399), .B1(n453), .Y(n196) );
  XOR2X1 U392 ( .A(b[13]), .B(n410), .Y(n452) );
  OAI22X1 U393 ( .A0(n453), .A1(n398), .B0(n399), .B1(n454), .Y(n195) );
  XOR2X1 U394 ( .A(b[14]), .B(n410), .Y(n453) );
  OAI22X1 U395 ( .A0(n454), .A1(n398), .B0(n399), .B1(n410), .Y(n194) );
  XOR2X1 U396 ( .A(b[15]), .B(n410), .Y(n454) );
  OAI2BB1X1 U397 ( .A0N(n398), .A1N(n399), .B0(a[3]), .Y(n193) );
  NOR2X1 U398 ( .A(n413), .B(n401), .Y(n192) );
  OAI22X1 U399 ( .A0(n456), .A1(n400), .B0(n401), .B1(n458), .Y(n191) );
  XOR2X1 U400 ( .A(n413), .B(a[5]), .Y(n456) );
  OAI22X1 U401 ( .A0(n458), .A1(n400), .B0(n401), .B1(n459), .Y(n190) );
  XOR2X1 U402 ( .A(b[1]), .B(n409), .Y(n458) );
  OAI22X1 U403 ( .A0(n459), .A1(n400), .B0(n401), .B1(n460), .Y(n189) );
  XOR2X1 U404 ( .A(b[2]), .B(n409), .Y(n459) );
  OAI22X1 U405 ( .A0(n460), .A1(n400), .B0(n401), .B1(n461), .Y(n188) );
  XOR2X1 U406 ( .A(b[3]), .B(n409), .Y(n460) );
  OAI22X1 U407 ( .A0(n461), .A1(n400), .B0(n401), .B1(n462), .Y(n187) );
  XOR2X1 U408 ( .A(b[4]), .B(n409), .Y(n461) );
  OAI22X1 U409 ( .A0(n462), .A1(n400), .B0(n401), .B1(n463), .Y(n186) );
  XOR2X1 U410 ( .A(b[5]), .B(n409), .Y(n462) );
  OAI22X1 U411 ( .A0(n463), .A1(n400), .B0(n401), .B1(n464), .Y(n185) );
  XOR2X1 U412 ( .A(b[6]), .B(n409), .Y(n463) );
  OAI22X1 U413 ( .A0(n464), .A1(n400), .B0(n401), .B1(n465), .Y(n184) );
  XOR2X1 U414 ( .A(b[7]), .B(n409), .Y(n464) );
  OAI22X1 U415 ( .A0(n465), .A1(n400), .B0(n401), .B1(n466), .Y(n183) );
  XOR2X1 U416 ( .A(b[8]), .B(n409), .Y(n465) );
  OAI22X1 U417 ( .A0(n466), .A1(n400), .B0(n401), .B1(n467), .Y(n182) );
  XOR2X1 U418 ( .A(b[9]), .B(n409), .Y(n466) );
  OAI22X1 U419 ( .A0(n467), .A1(n400), .B0(n401), .B1(n468), .Y(n181) );
  XOR2X1 U420 ( .A(b[10]), .B(n409), .Y(n467) );
  OAI22X1 U421 ( .A0(n468), .A1(n400), .B0(n401), .B1(n469), .Y(n180) );
  XOR2X1 U422 ( .A(b[11]), .B(n409), .Y(n468) );
  OAI22X1 U423 ( .A0(n469), .A1(n400), .B0(n401), .B1(n470), .Y(n179) );
  XOR2X1 U424 ( .A(b[12]), .B(n409), .Y(n469) );
  OAI22X1 U425 ( .A0(n470), .A1(n400), .B0(n401), .B1(n471), .Y(n178) );
  XOR2X1 U426 ( .A(b[13]), .B(n409), .Y(n470) );
  OAI22X1 U427 ( .A0(n471), .A1(n400), .B0(n401), .B1(n472), .Y(n177) );
  XOR2X1 U428 ( .A(b[14]), .B(n409), .Y(n471) );
  OAI22X1 U429 ( .A0(n472), .A1(n400), .B0(n401), .B1(n409), .Y(n176) );
  XOR2X1 U430 ( .A(b[15]), .B(n409), .Y(n472) );
  OAI2BB1X1 U431 ( .A0N(n400), .A1N(n401), .B0(a[5]), .Y(n175) );
  NOR2X1 U432 ( .A(n403), .B(n413), .Y(n174) );
  OAI22X1 U433 ( .A0(n473), .A1(n402), .B0(n403), .B1(n474), .Y(n173) );
  XOR2X1 U434 ( .A(n413), .B(n406), .Y(n473) );
  OAI22X1 U435 ( .A0(n474), .A1(n402), .B0(n403), .B1(n475), .Y(n172) );
  XOR2X1 U436 ( .A(b[1]), .B(n404), .Y(n474) );
  OAI22X1 U437 ( .A0(n475), .A1(n402), .B0(n403), .B1(n476), .Y(n171) );
  XOR2X1 U438 ( .A(b[2]), .B(n404), .Y(n475) );
  OAI22X1 U439 ( .A0(n476), .A1(n402), .B0(n403), .B1(n477), .Y(n170) );
  XOR2X1 U440 ( .A(b[3]), .B(n404), .Y(n476) );
  OAI22X1 U441 ( .A0(n477), .A1(n402), .B0(n403), .B1(n478), .Y(n169) );
  XOR2X1 U442 ( .A(b[4]), .B(n404), .Y(n477) );
  OAI22X1 U443 ( .A0(n478), .A1(n402), .B0(n403), .B1(n479), .Y(n168) );
  XOR2X1 U444 ( .A(b[5]), .B(n404), .Y(n478) );
  OAI22X1 U445 ( .A0(n479), .A1(n402), .B0(n403), .B1(n480), .Y(n167) );
  XOR2X1 U446 ( .A(b[6]), .B(n404), .Y(n479) );
  OAI22X1 U447 ( .A0(n480), .A1(n402), .B0(n403), .B1(n481), .Y(n166) );
  XOR2X1 U448 ( .A(b[7]), .B(n404), .Y(n480) );
  OAI22X1 U449 ( .A0(n481), .A1(n402), .B0(n403), .B1(n482), .Y(n165) );
  XOR2X1 U450 ( .A(b[8]), .B(n404), .Y(n481) );
  OAI22X1 U451 ( .A0(n482), .A1(n402), .B0(n403), .B1(n483), .Y(n164) );
  XOR2X1 U452 ( .A(b[9]), .B(n404), .Y(n482) );
  OAI22X1 U453 ( .A0(n483), .A1(n402), .B0(n403), .B1(n484), .Y(n163) );
  XOR2X1 U454 ( .A(b[10]), .B(n404), .Y(n483) );
  OAI22X1 U455 ( .A0(n484), .A1(n402), .B0(n403), .B1(n485), .Y(n162) );
  XOR2X1 U456 ( .A(b[11]), .B(n404), .Y(n484) );
  OAI22X1 U457 ( .A0(n485), .A1(n402), .B0(n403), .B1(n486), .Y(n161) );
  XOR2X1 U458 ( .A(b[12]), .B(n404), .Y(n485) );
  OAI22X1 U459 ( .A0(n486), .A1(n402), .B0(n403), .B1(n487), .Y(n160) );
  XOR2X1 U460 ( .A(b[13]), .B(n405), .Y(n486) );
  OAI22X1 U461 ( .A0(n487), .A1(n402), .B0(n403), .B1(n488), .Y(n159) );
  XOR2X1 U462 ( .A(b[14]), .B(n405), .Y(n487) );
  OAI22X1 U463 ( .A0(n488), .A1(n402), .B0(n403), .B1(n405), .Y(n158) );
  XOR2X1 U464 ( .A(b[15]), .B(n405), .Y(n488) );
  NOR2X1 U465 ( .A(n413), .B(n405), .Y(n156) );
  NOR2BX1 U466 ( .AN(b[1]), .B(n405), .Y(n155) );
  NOR2BX1 U467 ( .AN(b[2]), .B(n405), .Y(n154) );
  NOR2BX1 U468 ( .AN(b[3]), .B(n405), .Y(n153) );
  NOR2BX1 U469 ( .AN(b[4]), .B(n405), .Y(n152) );
  NOR2BX1 U470 ( .AN(b[5]), .B(n405), .Y(n151) );
  NOR2BX1 U471 ( .AN(b[6]), .B(n405), .Y(n150) );
  NOR2BX1 U472 ( .AN(b[7]), .B(n405), .Y(n149) );
  NOR2BX1 U473 ( .AN(b[8]), .B(n405), .Y(n148) );
  NOR2BX1 U474 ( .AN(b[10]), .B(n405), .Y(n147) );
  NOR2BX1 U475 ( .AN(b[11]), .B(n405), .Y(n146) );
  NOR2BX1 U476 ( .AN(b[13]), .B(n405), .Y(n145) );
  OAI21X1 U477 ( .A0(b[0]), .A1(n411), .B0(n397), .Y(n143) );
  OAI32XL U478 ( .A0(n410), .A1(b[0]), .A2(n399), .B0(n410), .B1(n398), .Y(
        n142) );
  XOR2X1 U479 ( .A(a[3]), .B(a[2]), .Y(n489) );
  OAI32XL U480 ( .A0(n409), .A1(b[0]), .A2(n401), .B0(n409), .B1(n400), .Y(
        n141) );
  XOR2X1 U481 ( .A(a[5]), .B(a[4]), .Y(n490) );
  OAI32XL U482 ( .A0(n405), .A1(b[0]), .A2(n403), .B0(n405), .B1(n402), .Y(
        n140) );
  XOR2X1 U483 ( .A(n406), .B(a[6]), .Y(n491) );
endmodule


module PE_1 ( pixel_00, pixel_01, pixel_02, pixel_10, pixel_11, pixel_12, 
        pixel_20, pixel_21, pixel_22, weight_00, weight_01, weight_02, 
        weight_10, weight_11, weight_12, weight_20, weight_21, weight_22, 
        out_pixel_00, out_pixel_01, out_pixel_02, out_pixel_10, out_pixel_11, 
        out_pixel_12, out_pixel_20, out_pixel_21, out_pixel_22, total, clk );
  input [7:0] pixel_00;
  input [7:0] pixel_01;
  input [7:0] pixel_02;
  input [7:0] pixel_10;
  input [7:0] pixel_11;
  input [7:0] pixel_12;
  input [7:0] pixel_20;
  input [7:0] pixel_21;
  input [7:0] pixel_22;
  input [15:0] weight_00;
  input [15:0] weight_01;
  input [15:0] weight_02;
  input [15:0] weight_10;
  input [15:0] weight_11;
  input [15:0] weight_12;
  input [15:0] weight_20;
  input [15:0] weight_21;
  input [15:0] weight_22;
  output [31:0] out_pixel_00;
  output [31:0] out_pixel_01;
  output [31:0] out_pixel_02;
  output [31:0] out_pixel_10;
  output [31:0] out_pixel_11;
  output [31:0] out_pixel_12;
  output [31:0] out_pixel_20;
  output [31:0] out_pixel_21;
  output [31:0] out_pixel_22;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, n1, n2, n3, n4, n5, n6, n7, n8,
         n9;
  assign out_pixel_00[31] = 1'b0;
  assign out_pixel_00[30] = 1'b0;
  assign out_pixel_00[29] = 1'b0;
  assign out_pixel_00[28] = 1'b0;
  assign out_pixel_00[27] = 1'b0;
  assign out_pixel_00[26] = 1'b0;
  assign out_pixel_00[25] = 1'b0;
  assign out_pixel_00[24] = 1'b0;
  assign out_pixel_01[31] = 1'b0;
  assign out_pixel_01[30] = 1'b0;
  assign out_pixel_01[29] = 1'b0;
  assign out_pixel_01[28] = 1'b0;
  assign out_pixel_01[27] = 1'b0;
  assign out_pixel_01[26] = 1'b0;
  assign out_pixel_01[25] = 1'b0;
  assign out_pixel_01[24] = 1'b0;
  assign out_pixel_02[31] = 1'b0;
  assign out_pixel_02[30] = 1'b0;
  assign out_pixel_02[29] = 1'b0;
  assign out_pixel_02[28] = 1'b0;
  assign out_pixel_02[27] = 1'b0;
  assign out_pixel_02[26] = 1'b0;
  assign out_pixel_02[25] = 1'b0;
  assign out_pixel_02[24] = 1'b0;
  assign out_pixel_10[31] = 1'b0;
  assign out_pixel_10[30] = 1'b0;
  assign out_pixel_10[29] = 1'b0;
  assign out_pixel_10[28] = 1'b0;
  assign out_pixel_10[27] = 1'b0;
  assign out_pixel_10[26] = 1'b0;
  assign out_pixel_10[25] = 1'b0;
  assign out_pixel_10[24] = 1'b0;
  assign out_pixel_11[31] = 1'b0;
  assign out_pixel_11[30] = 1'b0;
  assign out_pixel_11[29] = 1'b0;
  assign out_pixel_11[28] = 1'b0;
  assign out_pixel_11[27] = 1'b0;
  assign out_pixel_11[26] = 1'b0;
  assign out_pixel_11[25] = 1'b0;
  assign out_pixel_11[24] = 1'b0;
  assign out_pixel_12[31] = 1'b0;
  assign out_pixel_12[30] = 1'b0;
  assign out_pixel_12[29] = 1'b0;
  assign out_pixel_12[28] = 1'b0;
  assign out_pixel_12[27] = 1'b0;
  assign out_pixel_12[26] = 1'b0;
  assign out_pixel_12[25] = 1'b0;
  assign out_pixel_12[24] = 1'b0;
  assign out_pixel_20[31] = 1'b0;
  assign out_pixel_20[30] = 1'b0;
  assign out_pixel_20[29] = 1'b0;
  assign out_pixel_20[28] = 1'b0;
  assign out_pixel_20[27] = 1'b0;
  assign out_pixel_20[26] = 1'b0;
  assign out_pixel_20[25] = 1'b0;
  assign out_pixel_20[24] = 1'b0;
  assign out_pixel_21[31] = 1'b0;
  assign out_pixel_21[30] = 1'b0;
  assign out_pixel_21[29] = 1'b0;
  assign out_pixel_21[28] = 1'b0;
  assign out_pixel_21[27] = 1'b0;
  assign out_pixel_21[26] = 1'b0;
  assign out_pixel_21[25] = 1'b0;
  assign out_pixel_21[24] = 1'b0;
  assign out_pixel_22[31] = 1'b0;
  assign out_pixel_22[30] = 1'b0;
  assign out_pixel_22[29] = 1'b0;
  assign out_pixel_22[28] = 1'b0;
  assign out_pixel_22[27] = 1'b0;
  assign out_pixel_22[26] = 1'b0;
  assign out_pixel_22[25] = 1'b0;
  assign out_pixel_22[24] = 1'b0;

  PE_1_DW_mult_uns_8 mult_45 ( .a({n1, pixel_22[6:0]}), .b(weight_22), 
        .product({N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192}) );
  PE_1_DW_mult_uns_7 mult_44 ( .a({n2, pixel_21[6:0]}), .b(weight_21), 
        .product({N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, 
        N169, N168}) );
  PE_1_DW_mult_uns_6 mult_43 ( .a({n3, pixel_20[6:0]}), .b(weight_20), 
        .product({N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144}) );
  PE_1_DW_mult_uns_5 mult_42 ( .a({n4, pixel_12[6:0]}), .b(weight_12), 
        .product({N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}) );
  PE_1_DW_mult_uns_4 mult_41 ( .a({n5, pixel_11[6:0]}), .b(weight_11), 
        .product({N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96}) );
  PE_1_DW_mult_uns_3 mult_40 ( .a({n6, pixel_10[6:0]}), .b(weight_10), 
        .product({N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}) );
  PE_1_DW_mult_uns_2 mult_39 ( .a({n7, pixel_02[6:0]}), .b(weight_02), 
        .product({N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48}) );
  PE_1_DW_mult_uns_0 mult_38 ( .a({n8, pixel_01[6:0]}), .b(weight_01), 
        .product({N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24}) );
  PE_1_DW_mult_uns_1 mult_37 ( .a({n9, pixel_00[6:0]}), .b(weight_00), 
        .product({N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  DFFQXL \out_pixel_00_reg[23]  ( .D(N23), .CK(clk), .Q(out_pixel_00[23]) );
  DFFQXL \out_pixel_00_reg[22]  ( .D(N22), .CK(clk), .Q(out_pixel_00[22]) );
  DFFQXL \out_pixel_00_reg[21]  ( .D(N21), .CK(clk), .Q(out_pixel_00[21]) );
  DFFQXL \out_pixel_00_reg[20]  ( .D(N20), .CK(clk), .Q(out_pixel_00[20]) );
  DFFQXL \out_pixel_02_reg[23]  ( .D(N71), .CK(clk), .Q(out_pixel_02[23]) );
  DFFQXL \out_pixel_02_reg[22]  ( .D(N70), .CK(clk), .Q(out_pixel_02[22]) );
  DFFQXL \out_pixel_02_reg[21]  ( .D(N69), .CK(clk), .Q(out_pixel_02[21]) );
  DFFQXL \out_pixel_02_reg[20]  ( .D(N68), .CK(clk), .Q(out_pixel_02[20]) );
  DFFQXL \out_pixel_11_reg[23]  ( .D(N119), .CK(clk), .Q(out_pixel_11[23]) );
  DFFQXL \out_pixel_11_reg[22]  ( .D(N118), .CK(clk), .Q(out_pixel_11[22]) );
  DFFQXL \out_pixel_11_reg[21]  ( .D(N117), .CK(clk), .Q(out_pixel_11[21]) );
  DFFQXL \out_pixel_11_reg[20]  ( .D(N116), .CK(clk), .Q(out_pixel_11[20]) );
  DFFQXL \out_pixel_20_reg[23]  ( .D(N167), .CK(clk), .Q(out_pixel_20[23]) );
  DFFQXL \out_pixel_20_reg[22]  ( .D(N166), .CK(clk), .Q(out_pixel_20[22]) );
  DFFQXL \out_pixel_20_reg[21]  ( .D(N165), .CK(clk), .Q(out_pixel_20[21]) );
  DFFQXL \out_pixel_20_reg[20]  ( .D(N164), .CK(clk), .Q(out_pixel_20[20]) );
  DFFQXL \out_pixel_01_reg[23]  ( .D(N47), .CK(clk), .Q(out_pixel_01[23]) );
  DFFQXL \out_pixel_01_reg[22]  ( .D(N46), .CK(clk), .Q(out_pixel_01[22]) );
  DFFQXL \out_pixel_01_reg[21]  ( .D(N45), .CK(clk), .Q(out_pixel_01[21]) );
  DFFQXL \out_pixel_01_reg[20]  ( .D(N44), .CK(clk), .Q(out_pixel_01[20]) );
  DFFQXL \out_pixel_10_reg[23]  ( .D(N95), .CK(clk), .Q(out_pixel_10[23]) );
  DFFQXL \out_pixel_10_reg[22]  ( .D(N94), .CK(clk), .Q(out_pixel_10[22]) );
  DFFQXL \out_pixel_10_reg[21]  ( .D(N93), .CK(clk), .Q(out_pixel_10[21]) );
  DFFQXL \out_pixel_10_reg[20]  ( .D(N92), .CK(clk), .Q(out_pixel_10[20]) );
  DFFQXL \out_pixel_12_reg[23]  ( .D(N143), .CK(clk), .Q(out_pixel_12[23]) );
  DFFQXL \out_pixel_12_reg[22]  ( .D(N142), .CK(clk), .Q(out_pixel_12[22]) );
  DFFQXL \out_pixel_12_reg[21]  ( .D(N141), .CK(clk), .Q(out_pixel_12[21]) );
  DFFQXL \out_pixel_12_reg[20]  ( .D(N140), .CK(clk), .Q(out_pixel_12[20]) );
  DFFQXL \out_pixel_21_reg[23]  ( .D(N191), .CK(clk), .Q(out_pixel_21[23]) );
  DFFQXL \out_pixel_21_reg[22]  ( .D(N190), .CK(clk), .Q(out_pixel_21[22]) );
  DFFQXL \out_pixel_21_reg[21]  ( .D(N189), .CK(clk), .Q(out_pixel_21[21]) );
  DFFQXL \out_pixel_21_reg[20]  ( .D(N188), .CK(clk), .Q(out_pixel_21[20]) );
  DFFQXL \out_pixel_00_reg[19]  ( .D(N19), .CK(clk), .Q(out_pixel_00[19]) );
  DFFQXL \out_pixel_00_reg[18]  ( .D(N18), .CK(clk), .Q(out_pixel_00[18]) );
  DFFQXL \out_pixel_00_reg[17]  ( .D(N17), .CK(clk), .Q(out_pixel_00[17]) );
  DFFQXL \out_pixel_00_reg[16]  ( .D(N16), .CK(clk), .Q(out_pixel_00[16]) );
  DFFQXL \out_pixel_00_reg[15]  ( .D(N15), .CK(clk), .Q(out_pixel_00[15]) );
  DFFQXL \out_pixel_00_reg[14]  ( .D(N14), .CK(clk), .Q(out_pixel_00[14]) );
  DFFQXL \out_pixel_00_reg[13]  ( .D(N13), .CK(clk), .Q(out_pixel_00[13]) );
  DFFQXL \out_pixel_02_reg[19]  ( .D(N67), .CK(clk), .Q(out_pixel_02[19]) );
  DFFQXL \out_pixel_02_reg[18]  ( .D(N66), .CK(clk), .Q(out_pixel_02[18]) );
  DFFQXL \out_pixel_02_reg[17]  ( .D(N65), .CK(clk), .Q(out_pixel_02[17]) );
  DFFQXL \out_pixel_02_reg[16]  ( .D(N64), .CK(clk), .Q(out_pixel_02[16]) );
  DFFQXL \out_pixel_02_reg[15]  ( .D(N63), .CK(clk), .Q(out_pixel_02[15]) );
  DFFQXL \out_pixel_02_reg[14]  ( .D(N62), .CK(clk), .Q(out_pixel_02[14]) );
  DFFQXL \out_pixel_02_reg[13]  ( .D(N61), .CK(clk), .Q(out_pixel_02[13]) );
  DFFQXL \out_pixel_11_reg[19]  ( .D(N115), .CK(clk), .Q(out_pixel_11[19]) );
  DFFQXL \out_pixel_11_reg[18]  ( .D(N114), .CK(clk), .Q(out_pixel_11[18]) );
  DFFQXL \out_pixel_11_reg[17]  ( .D(N113), .CK(clk), .Q(out_pixel_11[17]) );
  DFFQXL \out_pixel_11_reg[16]  ( .D(N112), .CK(clk), .Q(out_pixel_11[16]) );
  DFFQXL \out_pixel_11_reg[15]  ( .D(N111), .CK(clk), .Q(out_pixel_11[15]) );
  DFFQXL \out_pixel_11_reg[14]  ( .D(N110), .CK(clk), .Q(out_pixel_11[14]) );
  DFFQXL \out_pixel_11_reg[13]  ( .D(N109), .CK(clk), .Q(out_pixel_11[13]) );
  DFFQXL \out_pixel_20_reg[19]  ( .D(N163), .CK(clk), .Q(out_pixel_20[19]) );
  DFFQXL \out_pixel_20_reg[18]  ( .D(N162), .CK(clk), .Q(out_pixel_20[18]) );
  DFFQXL \out_pixel_20_reg[17]  ( .D(N161), .CK(clk), .Q(out_pixel_20[17]) );
  DFFQXL \out_pixel_20_reg[16]  ( .D(N160), .CK(clk), .Q(out_pixel_20[16]) );
  DFFQXL \out_pixel_20_reg[15]  ( .D(N159), .CK(clk), .Q(out_pixel_20[15]) );
  DFFQXL \out_pixel_20_reg[14]  ( .D(N158), .CK(clk), .Q(out_pixel_20[14]) );
  DFFQXL \out_pixel_20_reg[13]  ( .D(N157), .CK(clk), .Q(out_pixel_20[13]) );
  DFFQXL \out_pixel_01_reg[19]  ( .D(N43), .CK(clk), .Q(out_pixel_01[19]) );
  DFFQXL \out_pixel_01_reg[18]  ( .D(N42), .CK(clk), .Q(out_pixel_01[18]) );
  DFFQXL \out_pixel_01_reg[17]  ( .D(N41), .CK(clk), .Q(out_pixel_01[17]) );
  DFFQXL \out_pixel_01_reg[16]  ( .D(N40), .CK(clk), .Q(out_pixel_01[16]) );
  DFFQXL \out_pixel_01_reg[15]  ( .D(N39), .CK(clk), .Q(out_pixel_01[15]) );
  DFFQXL \out_pixel_01_reg[14]  ( .D(N38), .CK(clk), .Q(out_pixel_01[14]) );
  DFFQXL \out_pixel_01_reg[13]  ( .D(N37), .CK(clk), .Q(out_pixel_01[13]) );
  DFFQXL \out_pixel_01_reg[12]  ( .D(N36), .CK(clk), .Q(out_pixel_01[12]) );
  DFFQXL \out_pixel_10_reg[19]  ( .D(N91), .CK(clk), .Q(out_pixel_10[19]) );
  DFFQXL \out_pixel_10_reg[18]  ( .D(N90), .CK(clk), .Q(out_pixel_10[18]) );
  DFFQXL \out_pixel_10_reg[17]  ( .D(N89), .CK(clk), .Q(out_pixel_10[17]) );
  DFFQXL \out_pixel_10_reg[16]  ( .D(N88), .CK(clk), .Q(out_pixel_10[16]) );
  DFFQXL \out_pixel_10_reg[15]  ( .D(N87), .CK(clk), .Q(out_pixel_10[15]) );
  DFFQXL \out_pixel_10_reg[14]  ( .D(N86), .CK(clk), .Q(out_pixel_10[14]) );
  DFFQXL \out_pixel_10_reg[13]  ( .D(N85), .CK(clk), .Q(out_pixel_10[13]) );
  DFFQXL \out_pixel_10_reg[12]  ( .D(N84), .CK(clk), .Q(out_pixel_10[12]) );
  DFFQXL \out_pixel_12_reg[19]  ( .D(N139), .CK(clk), .Q(out_pixel_12[19]) );
  DFFQXL \out_pixel_12_reg[18]  ( .D(N138), .CK(clk), .Q(out_pixel_12[18]) );
  DFFQXL \out_pixel_12_reg[17]  ( .D(N137), .CK(clk), .Q(out_pixel_12[17]) );
  DFFQXL \out_pixel_12_reg[16]  ( .D(N136), .CK(clk), .Q(out_pixel_12[16]) );
  DFFQXL \out_pixel_12_reg[15]  ( .D(N135), .CK(clk), .Q(out_pixel_12[15]) );
  DFFQXL \out_pixel_12_reg[14]  ( .D(N134), .CK(clk), .Q(out_pixel_12[14]) );
  DFFQXL \out_pixel_12_reg[13]  ( .D(N133), .CK(clk), .Q(out_pixel_12[13]) );
  DFFQXL \out_pixel_12_reg[12]  ( .D(N132), .CK(clk), .Q(out_pixel_12[12]) );
  DFFQXL \out_pixel_21_reg[19]  ( .D(N187), .CK(clk), .Q(out_pixel_21[19]) );
  DFFQXL \out_pixel_21_reg[18]  ( .D(N186), .CK(clk), .Q(out_pixel_21[18]) );
  DFFQXL \out_pixel_21_reg[17]  ( .D(N185), .CK(clk), .Q(out_pixel_21[17]) );
  DFFQXL \out_pixel_21_reg[16]  ( .D(N184), .CK(clk), .Q(out_pixel_21[16]) );
  DFFQXL \out_pixel_21_reg[15]  ( .D(N183), .CK(clk), .Q(out_pixel_21[15]) );
  DFFQXL \out_pixel_21_reg[14]  ( .D(N182), .CK(clk), .Q(out_pixel_21[14]) );
  DFFQXL \out_pixel_21_reg[13]  ( .D(N181), .CK(clk), .Q(out_pixel_21[13]) );
  DFFQXL \out_pixel_21_reg[12]  ( .D(N180), .CK(clk), .Q(out_pixel_21[12]) );
  DFFQXL \out_pixel_00_reg[12]  ( .D(N12), .CK(clk), .Q(out_pixel_00[12]) );
  DFFQXL \out_pixel_00_reg[11]  ( .D(N11), .CK(clk), .Q(out_pixel_00[11]) );
  DFFQXL \out_pixel_00_reg[10]  ( .D(N10), .CK(clk), .Q(out_pixel_00[10]) );
  DFFQXL \out_pixel_00_reg[9]  ( .D(N9), .CK(clk), .Q(out_pixel_00[9]) );
  DFFQXL \out_pixel_00_reg[8]  ( .D(N8), .CK(clk), .Q(out_pixel_00[8]) );
  DFFQXL \out_pixel_00_reg[7]  ( .D(N7), .CK(clk), .Q(out_pixel_00[7]) );
  DFFQXL \out_pixel_00_reg[6]  ( .D(N6), .CK(clk), .Q(out_pixel_00[6]) );
  DFFQXL \out_pixel_00_reg[5]  ( .D(N5), .CK(clk), .Q(out_pixel_00[5]) );
  DFFQXL \out_pixel_02_reg[12]  ( .D(N60), .CK(clk), .Q(out_pixel_02[12]) );
  DFFQXL \out_pixel_02_reg[11]  ( .D(N59), .CK(clk), .Q(out_pixel_02[11]) );
  DFFQXL \out_pixel_02_reg[10]  ( .D(N58), .CK(clk), .Q(out_pixel_02[10]) );
  DFFQXL \out_pixel_02_reg[9]  ( .D(N57), .CK(clk), .Q(out_pixel_02[9]) );
  DFFQXL \out_pixel_02_reg[8]  ( .D(N56), .CK(clk), .Q(out_pixel_02[8]) );
  DFFQXL \out_pixel_02_reg[7]  ( .D(N55), .CK(clk), .Q(out_pixel_02[7]) );
  DFFQXL \out_pixel_02_reg[6]  ( .D(N54), .CK(clk), .Q(out_pixel_02[6]) );
  DFFQXL \out_pixel_02_reg[5]  ( .D(N53), .CK(clk), .Q(out_pixel_02[5]) );
  DFFQXL \out_pixel_11_reg[12]  ( .D(N108), .CK(clk), .Q(out_pixel_11[12]) );
  DFFQXL \out_pixel_11_reg[11]  ( .D(N107), .CK(clk), .Q(out_pixel_11[11]) );
  DFFQXL \out_pixel_11_reg[10]  ( .D(N106), .CK(clk), .Q(out_pixel_11[10]) );
  DFFQXL \out_pixel_11_reg[9]  ( .D(N105), .CK(clk), .Q(out_pixel_11[9]) );
  DFFQXL \out_pixel_11_reg[8]  ( .D(N104), .CK(clk), .Q(out_pixel_11[8]) );
  DFFQXL \out_pixel_11_reg[7]  ( .D(N103), .CK(clk), .Q(out_pixel_11[7]) );
  DFFQXL \out_pixel_11_reg[6]  ( .D(N102), .CK(clk), .Q(out_pixel_11[6]) );
  DFFQXL \out_pixel_11_reg[5]  ( .D(N101), .CK(clk), .Q(out_pixel_11[5]) );
  DFFQXL \out_pixel_20_reg[12]  ( .D(N156), .CK(clk), .Q(out_pixel_20[12]) );
  DFFQXL \out_pixel_20_reg[11]  ( .D(N155), .CK(clk), .Q(out_pixel_20[11]) );
  DFFQXL \out_pixel_20_reg[10]  ( .D(N154), .CK(clk), .Q(out_pixel_20[10]) );
  DFFQXL \out_pixel_20_reg[9]  ( .D(N153), .CK(clk), .Q(out_pixel_20[9]) );
  DFFQXL \out_pixel_20_reg[8]  ( .D(N152), .CK(clk), .Q(out_pixel_20[8]) );
  DFFQXL \out_pixel_20_reg[7]  ( .D(N151), .CK(clk), .Q(out_pixel_20[7]) );
  DFFQXL \out_pixel_20_reg[6]  ( .D(N150), .CK(clk), .Q(out_pixel_20[6]) );
  DFFQXL \out_pixel_20_reg[5]  ( .D(N149), .CK(clk), .Q(out_pixel_20[5]) );
  DFFQXL \out_pixel_01_reg[11]  ( .D(N35), .CK(clk), .Q(out_pixel_01[11]) );
  DFFQXL \out_pixel_01_reg[10]  ( .D(N34), .CK(clk), .Q(out_pixel_01[10]) );
  DFFQXL \out_pixel_01_reg[9]  ( .D(N33), .CK(clk), .Q(out_pixel_01[9]) );
  DFFQXL \out_pixel_01_reg[8]  ( .D(N32), .CK(clk), .Q(out_pixel_01[8]) );
  DFFQXL \out_pixel_01_reg[7]  ( .D(N31), .CK(clk), .Q(out_pixel_01[7]) );
  DFFQXL \out_pixel_01_reg[6]  ( .D(N30), .CK(clk), .Q(out_pixel_01[6]) );
  DFFQXL \out_pixel_01_reg[5]  ( .D(N29), .CK(clk), .Q(out_pixel_01[5]) );
  DFFQXL \out_pixel_10_reg[11]  ( .D(N83), .CK(clk), .Q(out_pixel_10[11]) );
  DFFQXL \out_pixel_10_reg[10]  ( .D(N82), .CK(clk), .Q(out_pixel_10[10]) );
  DFFQXL \out_pixel_10_reg[9]  ( .D(N81), .CK(clk), .Q(out_pixel_10[9]) );
  DFFQXL \out_pixel_10_reg[8]  ( .D(N80), .CK(clk), .Q(out_pixel_10[8]) );
  DFFQXL \out_pixel_10_reg[7]  ( .D(N79), .CK(clk), .Q(out_pixel_10[7]) );
  DFFQXL \out_pixel_10_reg[6]  ( .D(N78), .CK(clk), .Q(out_pixel_10[6]) );
  DFFQXL \out_pixel_10_reg[5]  ( .D(N77), .CK(clk), .Q(out_pixel_10[5]) );
  DFFQXL \out_pixel_12_reg[11]  ( .D(N131), .CK(clk), .Q(out_pixel_12[11]) );
  DFFQXL \out_pixel_12_reg[10]  ( .D(N130), .CK(clk), .Q(out_pixel_12[10]) );
  DFFQXL \out_pixel_12_reg[9]  ( .D(N129), .CK(clk), .Q(out_pixel_12[9]) );
  DFFQXL \out_pixel_12_reg[8]  ( .D(N128), .CK(clk), .Q(out_pixel_12[8]) );
  DFFQXL \out_pixel_12_reg[7]  ( .D(N127), .CK(clk), .Q(out_pixel_12[7]) );
  DFFQXL \out_pixel_12_reg[6]  ( .D(N126), .CK(clk), .Q(out_pixel_12[6]) );
  DFFQXL \out_pixel_12_reg[5]  ( .D(N125), .CK(clk), .Q(out_pixel_12[5]) );
  DFFQXL \out_pixel_21_reg[11]  ( .D(N179), .CK(clk), .Q(out_pixel_21[11]) );
  DFFQXL \out_pixel_21_reg[10]  ( .D(N178), .CK(clk), .Q(out_pixel_21[10]) );
  DFFQXL \out_pixel_21_reg[9]  ( .D(N177), .CK(clk), .Q(out_pixel_21[9]) );
  DFFQXL \out_pixel_21_reg[8]  ( .D(N176), .CK(clk), .Q(out_pixel_21[8]) );
  DFFQXL \out_pixel_21_reg[7]  ( .D(N175), .CK(clk), .Q(out_pixel_21[7]) );
  DFFQXL \out_pixel_21_reg[6]  ( .D(N174), .CK(clk), .Q(out_pixel_21[6]) );
  DFFQXL \out_pixel_21_reg[5]  ( .D(N173), .CK(clk), .Q(out_pixel_21[5]) );
  DFFQXL \out_pixel_00_reg[4]  ( .D(N4), .CK(clk), .Q(out_pixel_00[4]) );
  DFFQXL \out_pixel_00_reg[3]  ( .D(N3), .CK(clk), .Q(out_pixel_00[3]) );
  DFFQXL \out_pixel_00_reg[2]  ( .D(N2), .CK(clk), .Q(out_pixel_00[2]) );
  DFFQXL \out_pixel_00_reg[1]  ( .D(N1), .CK(clk), .Q(out_pixel_00[1]) );
  DFFQXL \out_pixel_02_reg[4]  ( .D(N52), .CK(clk), .Q(out_pixel_02[4]) );
  DFFQXL \out_pixel_02_reg[3]  ( .D(N51), .CK(clk), .Q(out_pixel_02[3]) );
  DFFQXL \out_pixel_02_reg[2]  ( .D(N50), .CK(clk), .Q(out_pixel_02[2]) );
  DFFQXL \out_pixel_02_reg[1]  ( .D(N49), .CK(clk), .Q(out_pixel_02[1]) );
  DFFQXL \out_pixel_11_reg[4]  ( .D(N100), .CK(clk), .Q(out_pixel_11[4]) );
  DFFQXL \out_pixel_11_reg[3]  ( .D(N99), .CK(clk), .Q(out_pixel_11[3]) );
  DFFQXL \out_pixel_11_reg[2]  ( .D(N98), .CK(clk), .Q(out_pixel_11[2]) );
  DFFQXL \out_pixel_11_reg[1]  ( .D(N97), .CK(clk), .Q(out_pixel_11[1]) );
  DFFQXL \out_pixel_20_reg[4]  ( .D(N148), .CK(clk), .Q(out_pixel_20[4]) );
  DFFQXL \out_pixel_20_reg[3]  ( .D(N147), .CK(clk), .Q(out_pixel_20[3]) );
  DFFQXL \out_pixel_20_reg[2]  ( .D(N146), .CK(clk), .Q(out_pixel_20[2]) );
  DFFQXL \out_pixel_20_reg[1]  ( .D(N145), .CK(clk), .Q(out_pixel_20[1]) );
  DFFQXL \out_pixel_01_reg[4]  ( .D(N28), .CK(clk), .Q(out_pixel_01[4]) );
  DFFQXL \out_pixel_01_reg[3]  ( .D(N27), .CK(clk), .Q(out_pixel_01[3]) );
  DFFQXL \out_pixel_01_reg[2]  ( .D(N26), .CK(clk), .Q(out_pixel_01[2]) );
  DFFQXL \out_pixel_01_reg[1]  ( .D(N25), .CK(clk), .Q(out_pixel_01[1]) );
  DFFQXL \out_pixel_10_reg[4]  ( .D(N76), .CK(clk), .Q(out_pixel_10[4]) );
  DFFQXL \out_pixel_10_reg[3]  ( .D(N75), .CK(clk), .Q(out_pixel_10[3]) );
  DFFQXL \out_pixel_10_reg[2]  ( .D(N74), .CK(clk), .Q(out_pixel_10[2]) );
  DFFQXL \out_pixel_10_reg[1]  ( .D(N73), .CK(clk), .Q(out_pixel_10[1]) );
  DFFQXL \out_pixel_12_reg[4]  ( .D(N124), .CK(clk), .Q(out_pixel_12[4]) );
  DFFQXL \out_pixel_12_reg[3]  ( .D(N123), .CK(clk), .Q(out_pixel_12[3]) );
  DFFQXL \out_pixel_12_reg[2]  ( .D(N122), .CK(clk), .Q(out_pixel_12[2]) );
  DFFQXL \out_pixel_12_reg[1]  ( .D(N121), .CK(clk), .Q(out_pixel_12[1]) );
  DFFQXL \out_pixel_21_reg[4]  ( .D(N172), .CK(clk), .Q(out_pixel_21[4]) );
  DFFQXL \out_pixel_21_reg[3]  ( .D(N171), .CK(clk), .Q(out_pixel_21[3]) );
  DFFQXL \out_pixel_21_reg[2]  ( .D(N170), .CK(clk), .Q(out_pixel_21[2]) );
  DFFQXL \out_pixel_21_reg[1]  ( .D(N169), .CK(clk), .Q(out_pixel_21[1]) );
  DFFQXL \out_pixel_22_reg[23]  ( .D(N215), .CK(clk), .Q(out_pixel_22[23]) );
  DFFQXL \out_pixel_22_reg[3]  ( .D(N195), .CK(clk), .Q(out_pixel_22[3]) );
  DFFQXL \out_pixel_22_reg[1]  ( .D(N193), .CK(clk), .Q(out_pixel_22[1]) );
  DFFQXL \out_pixel_22_reg[22]  ( .D(N214), .CK(clk), .Q(out_pixel_22[22]) );
  DFFQXL \out_pixel_22_reg[21]  ( .D(N213), .CK(clk), .Q(out_pixel_22[21]) );
  DFFQXL \out_pixel_22_reg[6]  ( .D(N198), .CK(clk), .Q(out_pixel_22[6]) );
  DFFQXL \out_pixel_22_reg[5]  ( .D(N197), .CK(clk), .Q(out_pixel_22[5]) );
  DFFQXL \out_pixel_22_reg[4]  ( .D(N196), .CK(clk), .Q(out_pixel_22[4]) );
  DFFQXL \out_pixel_22_reg[2]  ( .D(N194), .CK(clk), .Q(out_pixel_22[2]) );
  DFFQXL \out_pixel_22_reg[0]  ( .D(N192), .CK(clk), .Q(out_pixel_22[0]) );
  DFFQXL \out_pixel_01_reg[0]  ( .D(N24), .CK(clk), .Q(out_pixel_01[0]) );
  DFFQXL \out_pixel_10_reg[0]  ( .D(N72), .CK(clk), .Q(out_pixel_10[0]) );
  DFFQXL \out_pixel_12_reg[0]  ( .D(N120), .CK(clk), .Q(out_pixel_12[0]) );
  DFFQXL \out_pixel_21_reg[0]  ( .D(N168), .CK(clk), .Q(out_pixel_21[0]) );
  DFFQXL \out_pixel_00_reg[0]  ( .D(N0), .CK(clk), .Q(out_pixel_00[0]) );
  DFFQXL \out_pixel_02_reg[0]  ( .D(N48), .CK(clk), .Q(out_pixel_02[0]) );
  DFFQXL \out_pixel_11_reg[0]  ( .D(N96), .CK(clk), .Q(out_pixel_11[0]) );
  DFFQXL \out_pixel_20_reg[0]  ( .D(N144), .CK(clk), .Q(out_pixel_20[0]) );
  DFFQXL \out_pixel_22_reg[20]  ( .D(N212), .CK(clk), .Q(out_pixel_22[20]) );
  DFFQXL \out_pixel_22_reg[19]  ( .D(N211), .CK(clk), .Q(out_pixel_22[19]) );
  DFFQXL \out_pixel_22_reg[18]  ( .D(N210), .CK(clk), .Q(out_pixel_22[18]) );
  DFFQXL \out_pixel_22_reg[17]  ( .D(N209), .CK(clk), .Q(out_pixel_22[17]) );
  DFFQXL \out_pixel_22_reg[16]  ( .D(N208), .CK(clk), .Q(out_pixel_22[16]) );
  DFFQXL \out_pixel_22_reg[15]  ( .D(N207), .CK(clk), .Q(out_pixel_22[15]) );
  DFFQXL \out_pixel_22_reg[14]  ( .D(N206), .CK(clk), .Q(out_pixel_22[14]) );
  DFFQXL \out_pixel_22_reg[13]  ( .D(N205), .CK(clk), .Q(out_pixel_22[13]) );
  DFFQXL \out_pixel_22_reg[12]  ( .D(N204), .CK(clk), .Q(out_pixel_22[12]) );
  DFFQXL \out_pixel_22_reg[11]  ( .D(N203), .CK(clk), .Q(out_pixel_22[11]) );
  DFFQXL \out_pixel_22_reg[10]  ( .D(N202), .CK(clk), .Q(out_pixel_22[10]) );
  DFFQXL \out_pixel_22_reg[9]  ( .D(N201), .CK(clk), .Q(out_pixel_22[9]) );
  DFFQXL \out_pixel_22_reg[8]  ( .D(N200), .CK(clk), .Q(out_pixel_22[8]) );
  DFFQXL \out_pixel_22_reg[7]  ( .D(N199), .CK(clk), .Q(out_pixel_22[7]) );
  BUFX2 U75 ( .A(pixel_22[7]), .Y(n1) );
  BUFX2 U76 ( .A(pixel_21[7]), .Y(n2) );
  BUFX2 U77 ( .A(pixel_20[7]), .Y(n3) );
  BUFX2 U78 ( .A(pixel_12[7]), .Y(n4) );
  BUFX2 U79 ( .A(pixel_11[7]), .Y(n5) );
  BUFX2 U80 ( .A(pixel_10[7]), .Y(n6) );
  BUFX2 U81 ( .A(pixel_02[7]), .Y(n7) );
  BUFX2 U82 ( .A(pixel_01[7]), .Y(n8) );
  BUFX2 U83 ( .A(pixel_00[7]), .Y(n9) );
endmodule


module Adder_tree_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_0 ( in1, in2, in3, in4, in5, in6, in7, in8, in9, total, clk
 );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  input [31:0] in5;
  input [31:0] in6;
  input [31:0] in7;
  input [31:0] in8;
  input [31:0] in9;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N223, N222, N221, N220, N219, N218, N217, N216,
         N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205,
         N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194,
         N193, N192;
  wire   [31:0] temp9;
  wire   [31:0] temp12;
  wire   [31:0] temp34;
  wire   [31:0] temp56;
  wire   [31:0] temp78;
  wire   [31:0] temp1234;
  wire   [31:0] temp5678;
  wire   [31:0] temp9_2;

  Adder_tree_0_DW01_add_0 add_29 ( .A(temp56), .B(temp78), .CI(1'b0), .SUM({
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160}) );
  Adder_tree_0_DW01_add_1 add_28 ( .A(temp12), .B(temp34), .CI(1'b0), .SUM({
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, 
        N135, N134, N133, N132, N131, N130, N129, N128}) );
  Adder_tree_0_DW01_add_2 add_25 ( .A(in7), .B(in8), .CI(1'b0), .SUM({N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96}) );
  Adder_tree_0_DW01_add_3 add_24 ( .A(in5), .B(in6), .CI(1'b0), .SUM({N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64}) );
  Adder_tree_0_DW01_add_4 add_23 ( .A(in3), .B(in4), .CI(1'b0), .SUM({N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32}) );
  Adder_tree_0_DW01_add_5 add_22 ( .A(in1), .B(in2), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Adder_tree_0_DW01_add_7 add_1_root_add_0_root_add_32_2 ( .A(temp9_2), .B(
        temp1234), .CI(1'b0), .SUM({N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 
        N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, 
        N192}) );
  Adder_tree_0_DW01_add_6 add_0_root_add_0_root_add_32_2 ( .A(temp5678), .B({
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192}), .CI(1'b0), .SUM({
        N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, 
        N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, 
        N231, N230, N229, N228, N227, N226, N225, N224}) );
  DFFQXL \temp9_2_reg[31]  ( .D(temp9[31]), .CK(clk), .Q(temp9_2[31]) );
  DFFQXL \temp9_2_reg[30]  ( .D(temp9[30]), .CK(clk), .Q(temp9_2[30]) );
  DFFQXL \temp9_2_reg[29]  ( .D(temp9[29]), .CK(clk), .Q(temp9_2[29]) );
  DFFQXL \temp12_reg[31]  ( .D(N31), .CK(clk), .Q(temp12[31]) );
  DFFQXL \temp12_reg[30]  ( .D(N30), .CK(clk), .Q(temp12[30]) );
  DFFQXL \temp12_reg[29]  ( .D(N29), .CK(clk), .Q(temp12[29]) );
  DFFQXL \temp12_reg[28]  ( .D(N28), .CK(clk), .Q(temp12[28]) );
  DFFQXL \temp12_reg[27]  ( .D(N27), .CK(clk), .Q(temp12[27]) );
  DFFQXL \temp56_reg[31]  ( .D(N95), .CK(clk), .Q(temp56[31]) );
  DFFQXL \temp56_reg[30]  ( .D(N94), .CK(clk), .Q(temp56[30]) );
  DFFQXL \temp56_reg[29]  ( .D(N93), .CK(clk), .Q(temp56[29]) );
  DFFQXL \temp56_reg[28]  ( .D(N92), .CK(clk), .Q(temp56[28]) );
  DFFQXL \temp56_reg[27]  ( .D(N91), .CK(clk), .Q(temp56[27]) );
  DFFQXL \temp5678_reg[31]  ( .D(N191), .CK(clk), .Q(temp5678[31]) );
  DFFQXL \temp5678_reg[30]  ( .D(N190), .CK(clk), .Q(temp5678[30]) );
  DFFQXL \temp5678_reg[29]  ( .D(N189), .CK(clk), .Q(temp5678[29]) );
  DFFQXL \temp5678_reg[28]  ( .D(N188), .CK(clk), .Q(temp5678[28]) );
  DFFQXL \temp5678_reg[27]  ( .D(N187), .CK(clk), .Q(temp5678[27]) );
  DFFQXL \temp34_reg[31]  ( .D(N63), .CK(clk), .Q(temp34[31]) );
  DFFQXL \temp34_reg[30]  ( .D(N62), .CK(clk), .Q(temp34[30]) );
  DFFQXL \temp34_reg[29]  ( .D(N61), .CK(clk), .Q(temp34[29]) );
  DFFQXL \temp34_reg[28]  ( .D(N60), .CK(clk), .Q(temp34[28]) );
  DFFQXL \temp34_reg[27]  ( .D(N59), .CK(clk), .Q(temp34[27]) );
  DFFQXL \temp78_reg[31]  ( .D(N127), .CK(clk), .Q(temp78[31]) );
  DFFQXL \temp78_reg[30]  ( .D(N126), .CK(clk), .Q(temp78[30]) );
  DFFQXL \temp78_reg[29]  ( .D(N125), .CK(clk), .Q(temp78[29]) );
  DFFQXL \temp78_reg[28]  ( .D(N124), .CK(clk), .Q(temp78[28]) );
  DFFQXL \temp78_reg[27]  ( .D(N123), .CK(clk), .Q(temp78[27]) );
  DFFQXL \temp1234_reg[31]  ( .D(N159), .CK(clk), .Q(temp1234[31]) );
  DFFQXL \temp1234_reg[30]  ( .D(N158), .CK(clk), .Q(temp1234[30]) );
  DFFQXL \temp1234_reg[29]  ( .D(N157), .CK(clk), .Q(temp1234[29]) );
  DFFQXL \temp9_2_reg[28]  ( .D(temp9[28]), .CK(clk), .Q(temp9_2[28]) );
  DFFQXL \temp9_2_reg[27]  ( .D(temp9[27]), .CK(clk), .Q(temp9_2[27]) );
  DFFQXL \temp9_2_reg[26]  ( .D(temp9[26]), .CK(clk), .Q(temp9_2[26]) );
  DFFQXL \temp9_2_reg[25]  ( .D(temp9[25]), .CK(clk), .Q(temp9_2[25]) );
  DFFQXL \temp9_2_reg[24]  ( .D(temp9[24]), .CK(clk), .Q(temp9_2[24]) );
  DFFQXL \temp9_2_reg[23]  ( .D(temp9[23]), .CK(clk), .Q(temp9_2[23]) );
  DFFQXL \temp9_2_reg[22]  ( .D(temp9[22]), .CK(clk), .Q(temp9_2[22]) );
  DFFQXL \temp12_reg[26]  ( .D(N26), .CK(clk), .Q(temp12[26]) );
  DFFQXL \temp12_reg[25]  ( .D(N25), .CK(clk), .Q(temp12[25]) );
  DFFQXL \temp12_reg[24]  ( .D(N24), .CK(clk), .Q(temp12[24]) );
  DFFQXL \temp12_reg[23]  ( .D(N23), .CK(clk), .Q(temp12[23]) );
  DFFQXL \temp12_reg[22]  ( .D(N22), .CK(clk), .Q(temp12[22]) );
  DFFQXL \temp12_reg[21]  ( .D(N21), .CK(clk), .Q(temp12[21]) );
  DFFQXL \temp12_reg[20]  ( .D(N20), .CK(clk), .Q(temp12[20]) );
  DFFQXL \temp56_reg[26]  ( .D(N90), .CK(clk), .Q(temp56[26]) );
  DFFQXL \temp56_reg[25]  ( .D(N89), .CK(clk), .Q(temp56[25]) );
  DFFQXL \temp56_reg[24]  ( .D(N88), .CK(clk), .Q(temp56[24]) );
  DFFQXL \temp56_reg[23]  ( .D(N87), .CK(clk), .Q(temp56[23]) );
  DFFQXL \temp56_reg[22]  ( .D(N86), .CK(clk), .Q(temp56[22]) );
  DFFQXL \temp56_reg[21]  ( .D(N85), .CK(clk), .Q(temp56[21]) );
  DFFQXL \temp56_reg[20]  ( .D(N84), .CK(clk), .Q(temp56[20]) );
  DFFQXL \temp5678_reg[26]  ( .D(N186), .CK(clk), .Q(temp5678[26]) );
  DFFQXL \temp5678_reg[25]  ( .D(N185), .CK(clk), .Q(temp5678[25]) );
  DFFQXL \temp5678_reg[24]  ( .D(N184), .CK(clk), .Q(temp5678[24]) );
  DFFQXL \temp5678_reg[23]  ( .D(N183), .CK(clk), .Q(temp5678[23]) );
  DFFQXL \temp5678_reg[22]  ( .D(N182), .CK(clk), .Q(temp5678[22]) );
  DFFQXL \temp5678_reg[21]  ( .D(N181), .CK(clk), .Q(temp5678[21]) );
  DFFQXL \temp5678_reg[20]  ( .D(N180), .CK(clk), .Q(temp5678[20]) );
  DFFQXL \temp34_reg[26]  ( .D(N58), .CK(clk), .Q(temp34[26]) );
  DFFQXL \temp34_reg[25]  ( .D(N57), .CK(clk), .Q(temp34[25]) );
  DFFQXL \temp34_reg[24]  ( .D(N56), .CK(clk), .Q(temp34[24]) );
  DFFQXL \temp34_reg[23]  ( .D(N55), .CK(clk), .Q(temp34[23]) );
  DFFQXL \temp34_reg[22]  ( .D(N54), .CK(clk), .Q(temp34[22]) );
  DFFQXL \temp34_reg[21]  ( .D(N53), .CK(clk), .Q(temp34[21]) );
  DFFQXL \temp34_reg[20]  ( .D(N52), .CK(clk), .Q(temp34[20]) );
  DFFQXL \temp78_reg[26]  ( .D(N122), .CK(clk), .Q(temp78[26]) );
  DFFQXL \temp78_reg[25]  ( .D(N121), .CK(clk), .Q(temp78[25]) );
  DFFQXL \temp78_reg[24]  ( .D(N120), .CK(clk), .Q(temp78[24]) );
  DFFQXL \temp78_reg[23]  ( .D(N119), .CK(clk), .Q(temp78[23]) );
  DFFQXL \temp78_reg[22]  ( .D(N118), .CK(clk), .Q(temp78[22]) );
  DFFQXL \temp78_reg[21]  ( .D(N117), .CK(clk), .Q(temp78[21]) );
  DFFQXL \temp78_reg[20]  ( .D(N116), .CK(clk), .Q(temp78[20]) );
  DFFQXL \temp1234_reg[28]  ( .D(N156), .CK(clk), .Q(temp1234[28]) );
  DFFQXL \temp1234_reg[27]  ( .D(N155), .CK(clk), .Q(temp1234[27]) );
  DFFQXL \temp1234_reg[26]  ( .D(N154), .CK(clk), .Q(temp1234[26]) );
  DFFQXL \temp1234_reg[25]  ( .D(N153), .CK(clk), .Q(temp1234[25]) );
  DFFQXL \temp1234_reg[24]  ( .D(N152), .CK(clk), .Q(temp1234[24]) );
  DFFQXL \temp1234_reg[23]  ( .D(N151), .CK(clk), .Q(temp1234[23]) );
  DFFQXL \temp1234_reg[22]  ( .D(N150), .CK(clk), .Q(temp1234[22]) );
  DFFQXL \temp1234_reg[21]  ( .D(N149), .CK(clk), .Q(temp1234[21]) );
  DFFQXL \temp9_2_reg[21]  ( .D(temp9[21]), .CK(clk), .Q(temp9_2[21]) );
  DFFQXL \temp9_2_reg[20]  ( .D(temp9[20]), .CK(clk), .Q(temp9_2[20]) );
  DFFQXL \temp9_2_reg[19]  ( .D(temp9[19]), .CK(clk), .Q(temp9_2[19]) );
  DFFQXL \temp9_2_reg[18]  ( .D(temp9[18]), .CK(clk), .Q(temp9_2[18]) );
  DFFQXL \temp9_2_reg[17]  ( .D(temp9[17]), .CK(clk), .Q(temp9_2[17]) );
  DFFQXL \temp9_2_reg[16]  ( .D(temp9[16]), .CK(clk), .Q(temp9_2[16]) );
  DFFQXL \temp9_2_reg[15]  ( .D(temp9[15]), .CK(clk), .Q(temp9_2[15]) );
  DFFQXL \temp9_2_reg[14]  ( .D(temp9[14]), .CK(clk), .Q(temp9_2[14]) );
  DFFQXL \temp12_reg[19]  ( .D(N19), .CK(clk), .Q(temp12[19]) );
  DFFQXL \temp12_reg[18]  ( .D(N18), .CK(clk), .Q(temp12[18]) );
  DFFQXL \temp12_reg[17]  ( .D(N17), .CK(clk), .Q(temp12[17]) );
  DFFQXL \temp12_reg[16]  ( .D(N16), .CK(clk), .Q(temp12[16]) );
  DFFQXL \temp12_reg[15]  ( .D(N15), .CK(clk), .Q(temp12[15]) );
  DFFQXL \temp12_reg[14]  ( .D(N14), .CK(clk), .Q(temp12[14]) );
  DFFQXL \temp12_reg[13]  ( .D(N13), .CK(clk), .Q(temp12[13]) );
  DFFQXL \temp12_reg[12]  ( .D(N12), .CK(clk), .Q(temp12[12]) );
  DFFQXL \temp56_reg[19]  ( .D(N83), .CK(clk), .Q(temp56[19]) );
  DFFQXL \temp56_reg[18]  ( .D(N82), .CK(clk), .Q(temp56[18]) );
  DFFQXL \temp56_reg[17]  ( .D(N81), .CK(clk), .Q(temp56[17]) );
  DFFQXL \temp56_reg[16]  ( .D(N80), .CK(clk), .Q(temp56[16]) );
  DFFQXL \temp56_reg[15]  ( .D(N79), .CK(clk), .Q(temp56[15]) );
  DFFQXL \temp56_reg[14]  ( .D(N78), .CK(clk), .Q(temp56[14]) );
  DFFQXL \temp56_reg[13]  ( .D(N77), .CK(clk), .Q(temp56[13]) );
  DFFQXL \temp56_reg[12]  ( .D(N76), .CK(clk), .Q(temp56[12]) );
  DFFQXL \temp5678_reg[19]  ( .D(N179), .CK(clk), .Q(temp5678[19]) );
  DFFQXL \temp5678_reg[18]  ( .D(N178), .CK(clk), .Q(temp5678[18]) );
  DFFQXL \temp5678_reg[17]  ( .D(N177), .CK(clk), .Q(temp5678[17]) );
  DFFQXL \temp5678_reg[16]  ( .D(N176), .CK(clk), .Q(temp5678[16]) );
  DFFQXL \temp5678_reg[15]  ( .D(N175), .CK(clk), .Q(temp5678[15]) );
  DFFQXL \temp5678_reg[14]  ( .D(N174), .CK(clk), .Q(temp5678[14]) );
  DFFQXL \temp5678_reg[13]  ( .D(N173), .CK(clk), .Q(temp5678[13]) );
  DFFQXL \temp5678_reg[12]  ( .D(N172), .CK(clk), .Q(temp5678[12]) );
  DFFQXL \temp34_reg[19]  ( .D(N51), .CK(clk), .Q(temp34[19]) );
  DFFQXL \temp34_reg[18]  ( .D(N50), .CK(clk), .Q(temp34[18]) );
  DFFQXL \temp34_reg[17]  ( .D(N49), .CK(clk), .Q(temp34[17]) );
  DFFQXL \temp34_reg[16]  ( .D(N48), .CK(clk), .Q(temp34[16]) );
  DFFQXL \temp34_reg[15]  ( .D(N47), .CK(clk), .Q(temp34[15]) );
  DFFQXL \temp34_reg[14]  ( .D(N46), .CK(clk), .Q(temp34[14]) );
  DFFQXL \temp34_reg[13]  ( .D(N45), .CK(clk), .Q(temp34[13]) );
  DFFQXL \temp34_reg[12]  ( .D(N44), .CK(clk), .Q(temp34[12]) );
  DFFQXL \temp78_reg[19]  ( .D(N115), .CK(clk), .Q(temp78[19]) );
  DFFQXL \temp78_reg[18]  ( .D(N114), .CK(clk), .Q(temp78[18]) );
  DFFQXL \temp78_reg[17]  ( .D(N113), .CK(clk), .Q(temp78[17]) );
  DFFQXL \temp78_reg[16]  ( .D(N112), .CK(clk), .Q(temp78[16]) );
  DFFQXL \temp78_reg[15]  ( .D(N111), .CK(clk), .Q(temp78[15]) );
  DFFQXL \temp78_reg[14]  ( .D(N110), .CK(clk), .Q(temp78[14]) );
  DFFQXL \temp78_reg[13]  ( .D(N109), .CK(clk), .Q(temp78[13]) );
  DFFQXL \temp78_reg[12]  ( .D(N108), .CK(clk), .Q(temp78[12]) );
  DFFQXL \temp1234_reg[20]  ( .D(N148), .CK(clk), .Q(temp1234[20]) );
  DFFQXL \temp1234_reg[19]  ( .D(N147), .CK(clk), .Q(temp1234[19]) );
  DFFQXL \temp1234_reg[18]  ( .D(N146), .CK(clk), .Q(temp1234[18]) );
  DFFQXL \temp1234_reg[17]  ( .D(N145), .CK(clk), .Q(temp1234[17]) );
  DFFQXL \temp1234_reg[16]  ( .D(N144), .CK(clk), .Q(temp1234[16]) );
  DFFQXL \temp1234_reg[15]  ( .D(N143), .CK(clk), .Q(temp1234[15]) );
  DFFQXL \temp1234_reg[14]  ( .D(N142), .CK(clk), .Q(temp1234[14]) );
  DFFQXL \temp9_2_reg[13]  ( .D(temp9[13]), .CK(clk), .Q(temp9_2[13]) );
  DFFQXL \temp9_2_reg[12]  ( .D(temp9[12]), .CK(clk), .Q(temp9_2[12]) );
  DFFQXL \temp9_2_reg[11]  ( .D(temp9[11]), .CK(clk), .Q(temp9_2[11]) );
  DFFQXL \temp9_2_reg[10]  ( .D(temp9[10]), .CK(clk), .Q(temp9_2[10]) );
  DFFQXL \temp9_2_reg[9]  ( .D(temp9[9]), .CK(clk), .Q(temp9_2[9]) );
  DFFQXL \temp9_2_reg[8]  ( .D(temp9[8]), .CK(clk), .Q(temp9_2[8]) );
  DFFQXL \temp9_2_reg[7]  ( .D(temp9[7]), .CK(clk), .Q(temp9_2[7]) );
  DFFQXL \temp12_reg[11]  ( .D(N11), .CK(clk), .Q(temp12[11]) );
  DFFQXL \temp12_reg[10]  ( .D(N10), .CK(clk), .Q(temp12[10]) );
  DFFQXL \temp12_reg[9]  ( .D(N9), .CK(clk), .Q(temp12[9]) );
  DFFQXL \temp12_reg[8]  ( .D(N8), .CK(clk), .Q(temp12[8]) );
  DFFQXL \temp12_reg[7]  ( .D(N7), .CK(clk), .Q(temp12[7]) );
  DFFQXL \temp12_reg[6]  ( .D(N6), .CK(clk), .Q(temp12[6]) );
  DFFQXL \temp12_reg[5]  ( .D(N5), .CK(clk), .Q(temp12[5]) );
  DFFQXL \temp56_reg[11]  ( .D(N75), .CK(clk), .Q(temp56[11]) );
  DFFQXL \temp56_reg[10]  ( .D(N74), .CK(clk), .Q(temp56[10]) );
  DFFQXL \temp56_reg[9]  ( .D(N73), .CK(clk), .Q(temp56[9]) );
  DFFQXL \temp56_reg[8]  ( .D(N72), .CK(clk), .Q(temp56[8]) );
  DFFQXL \temp56_reg[7]  ( .D(N71), .CK(clk), .Q(temp56[7]) );
  DFFQXL \temp56_reg[6]  ( .D(N70), .CK(clk), .Q(temp56[6]) );
  DFFQXL \temp56_reg[5]  ( .D(N69), .CK(clk), .Q(temp56[5]) );
  DFFQXL \temp5678_reg[11]  ( .D(N171), .CK(clk), .Q(temp5678[11]) );
  DFFQXL \temp5678_reg[10]  ( .D(N170), .CK(clk), .Q(temp5678[10]) );
  DFFQXL \temp5678_reg[9]  ( .D(N169), .CK(clk), .Q(temp5678[9]) );
  DFFQXL \temp5678_reg[8]  ( .D(N168), .CK(clk), .Q(temp5678[8]) );
  DFFQXL \temp5678_reg[7]  ( .D(N167), .CK(clk), .Q(temp5678[7]) );
  DFFQXL \temp5678_reg[6]  ( .D(N166), .CK(clk), .Q(temp5678[6]) );
  DFFQXL \temp5678_reg[5]  ( .D(N165), .CK(clk), .Q(temp5678[5]) );
  DFFQXL \temp34_reg[11]  ( .D(N43), .CK(clk), .Q(temp34[11]) );
  DFFQXL \temp34_reg[10]  ( .D(N42), .CK(clk), .Q(temp34[10]) );
  DFFQXL \temp34_reg[9]  ( .D(N41), .CK(clk), .Q(temp34[9]) );
  DFFQXL \temp34_reg[8]  ( .D(N40), .CK(clk), .Q(temp34[8]) );
  DFFQXL \temp34_reg[7]  ( .D(N39), .CK(clk), .Q(temp34[7]) );
  DFFQXL \temp34_reg[6]  ( .D(N38), .CK(clk), .Q(temp34[6]) );
  DFFQXL \temp34_reg[5]  ( .D(N37), .CK(clk), .Q(temp34[5]) );
  DFFQXL \temp78_reg[11]  ( .D(N107), .CK(clk), .Q(temp78[11]) );
  DFFQXL \temp78_reg[10]  ( .D(N106), .CK(clk), .Q(temp78[10]) );
  DFFQXL \temp78_reg[9]  ( .D(N105), .CK(clk), .Q(temp78[9]) );
  DFFQXL \temp78_reg[8]  ( .D(N104), .CK(clk), .Q(temp78[8]) );
  DFFQXL \temp78_reg[7]  ( .D(N103), .CK(clk), .Q(temp78[7]) );
  DFFQXL \temp78_reg[6]  ( .D(N102), .CK(clk), .Q(temp78[6]) );
  DFFQXL \temp78_reg[5]  ( .D(N101), .CK(clk), .Q(temp78[5]) );
  DFFQXL \temp1234_reg[13]  ( .D(N141), .CK(clk), .Q(temp1234[13]) );
  DFFQXL \temp1234_reg[12]  ( .D(N140), .CK(clk), .Q(temp1234[12]) );
  DFFQXL \temp1234_reg[11]  ( .D(N139), .CK(clk), .Q(temp1234[11]) );
  DFFQXL \temp1234_reg[10]  ( .D(N138), .CK(clk), .Q(temp1234[10]) );
  DFFQXL \temp1234_reg[9]  ( .D(N137), .CK(clk), .Q(temp1234[9]) );
  DFFQXL \temp1234_reg[8]  ( .D(N136), .CK(clk), .Q(temp1234[8]) );
  DFFQXL \temp1234_reg[7]  ( .D(N135), .CK(clk), .Q(temp1234[7]) );
  DFFQXL \temp1234_reg[6]  ( .D(N134), .CK(clk), .Q(temp1234[6]) );
  DFFQXL \temp9_2_reg[6]  ( .D(temp9[6]), .CK(clk), .Q(temp9_2[6]) );
  DFFQXL \temp9_2_reg[5]  ( .D(temp9[5]), .CK(clk), .Q(temp9_2[5]) );
  DFFQXL \temp9_2_reg[4]  ( .D(temp9[4]), .CK(clk), .Q(temp9_2[4]) );
  DFFQXL \temp9_2_reg[3]  ( .D(temp9[3]), .CK(clk), .Q(temp9_2[3]) );
  DFFQXL \temp9_2_reg[2]  ( .D(temp9[2]), .CK(clk), .Q(temp9_2[2]) );
  DFFQXL \temp9_2_reg[1]  ( .D(temp9[1]), .CK(clk), .Q(temp9_2[1]) );
  DFFQXL \temp12_reg[4]  ( .D(N4), .CK(clk), .Q(temp12[4]) );
  DFFQXL \temp12_reg[3]  ( .D(N3), .CK(clk), .Q(temp12[3]) );
  DFFQXL \temp12_reg[2]  ( .D(N2), .CK(clk), .Q(temp12[2]) );
  DFFQXL \temp12_reg[1]  ( .D(N1), .CK(clk), .Q(temp12[1]) );
  DFFQXL \temp56_reg[4]  ( .D(N68), .CK(clk), .Q(temp56[4]) );
  DFFQXL \temp56_reg[3]  ( .D(N67), .CK(clk), .Q(temp56[3]) );
  DFFQXL \temp56_reg[2]  ( .D(N66), .CK(clk), .Q(temp56[2]) );
  DFFQXL \temp56_reg[1]  ( .D(N65), .CK(clk), .Q(temp56[1]) );
  DFFQXL \temp5678_reg[4]  ( .D(N164), .CK(clk), .Q(temp5678[4]) );
  DFFQXL \temp5678_reg[3]  ( .D(N163), .CK(clk), .Q(temp5678[3]) );
  DFFQXL \temp5678_reg[2]  ( .D(N162), .CK(clk), .Q(temp5678[2]) );
  DFFQXL \temp5678_reg[1]  ( .D(N161), .CK(clk), .Q(temp5678[1]) );
  DFFQXL \temp34_reg[4]  ( .D(N36), .CK(clk), .Q(temp34[4]) );
  DFFQXL \temp34_reg[3]  ( .D(N35), .CK(clk), .Q(temp34[3]) );
  DFFQXL \temp34_reg[2]  ( .D(N34), .CK(clk), .Q(temp34[2]) );
  DFFQXL \temp34_reg[1]  ( .D(N33), .CK(clk), .Q(temp34[1]) );
  DFFQXL \temp78_reg[4]  ( .D(N100), .CK(clk), .Q(temp78[4]) );
  DFFQXL \temp78_reg[3]  ( .D(N99), .CK(clk), .Q(temp78[3]) );
  DFFQXL \temp78_reg[2]  ( .D(N98), .CK(clk), .Q(temp78[2]) );
  DFFQXL \temp78_reg[1]  ( .D(N97), .CK(clk), .Q(temp78[1]) );
  DFFQXL \temp1234_reg[5]  ( .D(N133), .CK(clk), .Q(temp1234[5]) );
  DFFQXL \temp1234_reg[4]  ( .D(N132), .CK(clk), .Q(temp1234[4]) );
  DFFQXL \temp1234_reg[3]  ( .D(N131), .CK(clk), .Q(temp1234[3]) );
  DFFQXL \temp1234_reg[2]  ( .D(N130), .CK(clk), .Q(temp1234[2]) );
  DFFQXL \temp1234_reg[1]  ( .D(N129), .CK(clk), .Q(temp1234[1]) );
  DFFQXL \total_reg[31]  ( .D(N255), .CK(clk), .Q(total[31]) );
  DFFQXL \total_reg[30]  ( .D(N254), .CK(clk), .Q(total[30]) );
  DFFQXL \total_reg[29]  ( .D(N253), .CK(clk), .Q(total[29]) );
  DFFQXL \total_reg[28]  ( .D(N252), .CK(clk), .Q(total[28]) );
  DFFQXL \total_reg[27]  ( .D(N251), .CK(clk), .Q(total[27]) );
  DFFQXL \total_reg[26]  ( .D(N250), .CK(clk), .Q(total[26]) );
  DFFQXL \total_reg[25]  ( .D(N249), .CK(clk), .Q(total[25]) );
  DFFQXL \total_reg[24]  ( .D(N248), .CK(clk), .Q(total[24]) );
  DFFQXL \total_reg[23]  ( .D(N247), .CK(clk), .Q(total[23]) );
  DFFQXL \total_reg[22]  ( .D(N246), .CK(clk), .Q(total[22]) );
  DFFQXL \total_reg[21]  ( .D(N245), .CK(clk), .Q(total[21]) );
  DFFQXL \total_reg[20]  ( .D(N244), .CK(clk), .Q(total[20]) );
  DFFQXL \total_reg[19]  ( .D(N243), .CK(clk), .Q(total[19]) );
  DFFQXL \total_reg[18]  ( .D(N242), .CK(clk), .Q(total[18]) );
  DFFQXL \total_reg[17]  ( .D(N241), .CK(clk), .Q(total[17]) );
  DFFQXL \total_reg[16]  ( .D(N240), .CK(clk), .Q(total[16]) );
  DFFQXL \total_reg[15]  ( .D(N239), .CK(clk), .Q(total[15]) );
  DFFQXL \total_reg[14]  ( .D(N238), .CK(clk), .Q(total[14]) );
  DFFQXL \total_reg[13]  ( .D(N237), .CK(clk), .Q(total[13]) );
  DFFQXL \total_reg[12]  ( .D(N236), .CK(clk), .Q(total[12]) );
  DFFQXL \total_reg[11]  ( .D(N235), .CK(clk), .Q(total[11]) );
  DFFQXL \total_reg[10]  ( .D(N234), .CK(clk), .Q(total[10]) );
  DFFQXL \total_reg[9]  ( .D(N233), .CK(clk), .Q(total[9]) );
  DFFQXL \total_reg[8]  ( .D(N232), .CK(clk), .Q(total[8]) );
  DFFQXL \total_reg[7]  ( .D(N231), .CK(clk), .Q(total[7]) );
  DFFQXL \total_reg[6]  ( .D(N230), .CK(clk), .Q(total[6]) );
  DFFQXL \total_reg[5]  ( .D(N229), .CK(clk), .Q(total[5]) );
  DFFQXL \total_reg[4]  ( .D(N228), .CK(clk), .Q(total[4]) );
  DFFQXL \total_reg[3]  ( .D(N227), .CK(clk), .Q(total[3]) );
  DFFQXL \total_reg[2]  ( .D(N226), .CK(clk), .Q(total[2]) );
  DFFQXL \total_reg[1]  ( .D(N225), .CK(clk), .Q(total[1]) );
  DFFQXL \total_reg[0]  ( .D(N224), .CK(clk), .Q(total[0]) );
  DFFQXL \temp34_reg[0]  ( .D(N32), .CK(clk), .Q(temp34[0]) );
  DFFQXL \temp78_reg[0]  ( .D(N96), .CK(clk), .Q(temp78[0]) );
  DFFQXL \temp1234_reg[0]  ( .D(N128), .CK(clk), .Q(temp1234[0]) );
  DFFQXL \temp12_reg[0]  ( .D(N0), .CK(clk), .Q(temp12[0]) );
  DFFQXL \temp56_reg[0]  ( .D(N64), .CK(clk), .Q(temp56[0]) );
  DFFQXL \temp5678_reg[0]  ( .D(N160), .CK(clk), .Q(temp5678[0]) );
  DFFQXL \temp9_2_reg[0]  ( .D(temp9[0]), .CK(clk), .Q(temp9_2[0]) );
  DFFQXL \temp9_reg[31]  ( .D(in9[31]), .CK(clk), .Q(temp9[31]) );
  DFFQXL \temp9_reg[30]  ( .D(in9[30]), .CK(clk), .Q(temp9[30]) );
  DFFQXL \temp9_reg[29]  ( .D(in9[29]), .CK(clk), .Q(temp9[29]) );
  DFFQXL \temp9_reg[28]  ( .D(in9[28]), .CK(clk), .Q(temp9[28]) );
  DFFQXL \temp9_reg[27]  ( .D(in9[27]), .CK(clk), .Q(temp9[27]) );
  DFFQXL \temp9_reg[26]  ( .D(in9[26]), .CK(clk), .Q(temp9[26]) );
  DFFQXL \temp9_reg[25]  ( .D(in9[25]), .CK(clk), .Q(temp9[25]) );
  DFFQXL \temp9_reg[24]  ( .D(in9[24]), .CK(clk), .Q(temp9[24]) );
  DFFQXL \temp9_reg[23]  ( .D(in9[23]), .CK(clk), .Q(temp9[23]) );
  DFFQXL \temp9_reg[22]  ( .D(in9[22]), .CK(clk), .Q(temp9[22]) );
  DFFQXL \temp9_reg[21]  ( .D(in9[21]), .CK(clk), .Q(temp9[21]) );
  DFFQXL \temp9_reg[20]  ( .D(in9[20]), .CK(clk), .Q(temp9[20]) );
  DFFQXL \temp9_reg[19]  ( .D(in9[19]), .CK(clk), .Q(temp9[19]) );
  DFFQXL \temp9_reg[18]  ( .D(in9[18]), .CK(clk), .Q(temp9[18]) );
  DFFQXL \temp9_reg[17]  ( .D(in9[17]), .CK(clk), .Q(temp9[17]) );
  DFFQXL \temp9_reg[16]  ( .D(in9[16]), .CK(clk), .Q(temp9[16]) );
  DFFQXL \temp9_reg[15]  ( .D(in9[15]), .CK(clk), .Q(temp9[15]) );
  DFFQXL \temp9_reg[14]  ( .D(in9[14]), .CK(clk), .Q(temp9[14]) );
  DFFQXL \temp9_reg[13]  ( .D(in9[13]), .CK(clk), .Q(temp9[13]) );
  DFFQXL \temp9_reg[12]  ( .D(in9[12]), .CK(clk), .Q(temp9[12]) );
  DFFQXL \temp9_reg[11]  ( .D(in9[11]), .CK(clk), .Q(temp9[11]) );
  DFFQXL \temp9_reg[10]  ( .D(in9[10]), .CK(clk), .Q(temp9[10]) );
  DFFQXL \temp9_reg[9]  ( .D(in9[9]), .CK(clk), .Q(temp9[9]) );
  DFFQXL \temp9_reg[8]  ( .D(in9[8]), .CK(clk), .Q(temp9[8]) );
  DFFQXL \temp9_reg[7]  ( .D(in9[7]), .CK(clk), .Q(temp9[7]) );
  DFFQXL \temp9_reg[6]  ( .D(in9[6]), .CK(clk), .Q(temp9[6]) );
  DFFQXL \temp9_reg[5]  ( .D(in9[5]), .CK(clk), .Q(temp9[5]) );
  DFFQXL \temp9_reg[4]  ( .D(in9[4]), .CK(clk), .Q(temp9[4]) );
  DFFQXL \temp9_reg[3]  ( .D(in9[3]), .CK(clk), .Q(temp9[3]) );
  DFFQXL \temp9_reg[2]  ( .D(in9[2]), .CK(clk), .Q(temp9[2]) );
  DFFQXL \temp9_reg[1]  ( .D(in9[1]), .CK(clk), .Q(temp9[1]) );
  DFFQXL \temp9_reg[0]  ( .D(in9[0]), .CK(clk), .Q(temp9[0]) );
endmodule


module Adder_tree_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_3 ( in1, in2, in3, in4, in5, in6, in7, in8, in9, total, clk
 );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  input [31:0] in5;
  input [31:0] in6;
  input [31:0] in7;
  input [31:0] in8;
  input [31:0] in9;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N223, N222, N221, N220, N219, N218, N217, N216,
         N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205,
         N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194,
         N193, N192;
  wire   [31:0] temp9;
  wire   [31:0] temp12;
  wire   [31:0] temp34;
  wire   [31:0] temp56;
  wire   [31:0] temp78;
  wire   [31:0] temp1234;
  wire   [31:0] temp5678;
  wire   [31:0] temp9_2;

  Adder_tree_3_DW01_add_0 add_29 ( .A(temp56), .B(temp78), .CI(1'b0), .SUM({
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160}) );
  Adder_tree_3_DW01_add_1 add_28 ( .A(temp12), .B(temp34), .CI(1'b0), .SUM({
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, 
        N135, N134, N133, N132, N131, N130, N129, N128}) );
  Adder_tree_3_DW01_add_2 add_25 ( .A(in7), .B(in8), .CI(1'b0), .SUM({N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96}) );
  Adder_tree_3_DW01_add_3 add_24 ( .A(in5), .B(in6), .CI(1'b0), .SUM({N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64}) );
  Adder_tree_3_DW01_add_4 add_23 ( .A(in3), .B(in4), .CI(1'b0), .SUM({N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32}) );
  Adder_tree_3_DW01_add_5 add_22 ( .A(in1), .B(in2), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Adder_tree_3_DW01_add_7 add_1_root_add_0_root_add_32_2 ( .A(temp9_2), .B(
        temp1234), .CI(1'b0), .SUM({N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 
        N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, 
        N192}) );
  Adder_tree_3_DW01_add_6 add_0_root_add_0_root_add_32_2 ( .A(temp5678), .B({
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192}), .CI(1'b0), .SUM({
        N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, 
        N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, 
        N231, N230, N229, N228, N227, N226, N225, N224}) );
  DFFQXL \temp9_2_reg[31]  ( .D(temp9[31]), .CK(clk), .Q(temp9_2[31]) );
  DFFQXL \temp9_2_reg[30]  ( .D(temp9[30]), .CK(clk), .Q(temp9_2[30]) );
  DFFQXL \temp9_2_reg[29]  ( .D(temp9[29]), .CK(clk), .Q(temp9_2[29]) );
  DFFQXL \temp12_reg[31]  ( .D(N31), .CK(clk), .Q(temp12[31]) );
  DFFQXL \temp12_reg[30]  ( .D(N30), .CK(clk), .Q(temp12[30]) );
  DFFQXL \temp12_reg[29]  ( .D(N29), .CK(clk), .Q(temp12[29]) );
  DFFQXL \temp12_reg[28]  ( .D(N28), .CK(clk), .Q(temp12[28]) );
  DFFQXL \temp12_reg[27]  ( .D(N27), .CK(clk), .Q(temp12[27]) );
  DFFQXL \temp56_reg[31]  ( .D(N95), .CK(clk), .Q(temp56[31]) );
  DFFQXL \temp56_reg[30]  ( .D(N94), .CK(clk), .Q(temp56[30]) );
  DFFQXL \temp56_reg[29]  ( .D(N93), .CK(clk), .Q(temp56[29]) );
  DFFQXL \temp56_reg[28]  ( .D(N92), .CK(clk), .Q(temp56[28]) );
  DFFQXL \temp56_reg[27]  ( .D(N91), .CK(clk), .Q(temp56[27]) );
  DFFQXL \temp5678_reg[31]  ( .D(N191), .CK(clk), .Q(temp5678[31]) );
  DFFQXL \temp5678_reg[30]  ( .D(N190), .CK(clk), .Q(temp5678[30]) );
  DFFQXL \temp5678_reg[29]  ( .D(N189), .CK(clk), .Q(temp5678[29]) );
  DFFQXL \temp5678_reg[28]  ( .D(N188), .CK(clk), .Q(temp5678[28]) );
  DFFQXL \temp5678_reg[27]  ( .D(N187), .CK(clk), .Q(temp5678[27]) );
  DFFQXL \temp34_reg[31]  ( .D(N63), .CK(clk), .Q(temp34[31]) );
  DFFQXL \temp34_reg[30]  ( .D(N62), .CK(clk), .Q(temp34[30]) );
  DFFQXL \temp34_reg[29]  ( .D(N61), .CK(clk), .Q(temp34[29]) );
  DFFQXL \temp34_reg[28]  ( .D(N60), .CK(clk), .Q(temp34[28]) );
  DFFQXL \temp34_reg[27]  ( .D(N59), .CK(clk), .Q(temp34[27]) );
  DFFQXL \temp78_reg[31]  ( .D(N127), .CK(clk), .Q(temp78[31]) );
  DFFQXL \temp78_reg[30]  ( .D(N126), .CK(clk), .Q(temp78[30]) );
  DFFQXL \temp78_reg[29]  ( .D(N125), .CK(clk), .Q(temp78[29]) );
  DFFQXL \temp78_reg[28]  ( .D(N124), .CK(clk), .Q(temp78[28]) );
  DFFQXL \temp78_reg[27]  ( .D(N123), .CK(clk), .Q(temp78[27]) );
  DFFQXL \temp1234_reg[31]  ( .D(N159), .CK(clk), .Q(temp1234[31]) );
  DFFQXL \temp1234_reg[30]  ( .D(N158), .CK(clk), .Q(temp1234[30]) );
  DFFQXL \temp1234_reg[29]  ( .D(N157), .CK(clk), .Q(temp1234[29]) );
  DFFQXL \temp9_2_reg[28]  ( .D(temp9[28]), .CK(clk), .Q(temp9_2[28]) );
  DFFQXL \temp9_2_reg[27]  ( .D(temp9[27]), .CK(clk), .Q(temp9_2[27]) );
  DFFQXL \temp9_2_reg[26]  ( .D(temp9[26]), .CK(clk), .Q(temp9_2[26]) );
  DFFQXL \temp9_2_reg[25]  ( .D(temp9[25]), .CK(clk), .Q(temp9_2[25]) );
  DFFQXL \temp9_2_reg[24]  ( .D(temp9[24]), .CK(clk), .Q(temp9_2[24]) );
  DFFQXL \temp9_2_reg[23]  ( .D(temp9[23]), .CK(clk), .Q(temp9_2[23]) );
  DFFQXL \temp9_2_reg[22]  ( .D(temp9[22]), .CK(clk), .Q(temp9_2[22]) );
  DFFQXL \temp12_reg[26]  ( .D(N26), .CK(clk), .Q(temp12[26]) );
  DFFQXL \temp12_reg[25]  ( .D(N25), .CK(clk), .Q(temp12[25]) );
  DFFQXL \temp12_reg[24]  ( .D(N24), .CK(clk), .Q(temp12[24]) );
  DFFQXL \temp12_reg[23]  ( .D(N23), .CK(clk), .Q(temp12[23]) );
  DFFQXL \temp12_reg[22]  ( .D(N22), .CK(clk), .Q(temp12[22]) );
  DFFQXL \temp12_reg[21]  ( .D(N21), .CK(clk), .Q(temp12[21]) );
  DFFQXL \temp12_reg[20]  ( .D(N20), .CK(clk), .Q(temp12[20]) );
  DFFQXL \temp56_reg[26]  ( .D(N90), .CK(clk), .Q(temp56[26]) );
  DFFQXL \temp56_reg[25]  ( .D(N89), .CK(clk), .Q(temp56[25]) );
  DFFQXL \temp56_reg[24]  ( .D(N88), .CK(clk), .Q(temp56[24]) );
  DFFQXL \temp56_reg[23]  ( .D(N87), .CK(clk), .Q(temp56[23]) );
  DFFQXL \temp56_reg[22]  ( .D(N86), .CK(clk), .Q(temp56[22]) );
  DFFQXL \temp56_reg[21]  ( .D(N85), .CK(clk), .Q(temp56[21]) );
  DFFQXL \temp56_reg[20]  ( .D(N84), .CK(clk), .Q(temp56[20]) );
  DFFQXL \temp5678_reg[26]  ( .D(N186), .CK(clk), .Q(temp5678[26]) );
  DFFQXL \temp5678_reg[25]  ( .D(N185), .CK(clk), .Q(temp5678[25]) );
  DFFQXL \temp5678_reg[24]  ( .D(N184), .CK(clk), .Q(temp5678[24]) );
  DFFQXL \temp5678_reg[23]  ( .D(N183), .CK(clk), .Q(temp5678[23]) );
  DFFQXL \temp5678_reg[22]  ( .D(N182), .CK(clk), .Q(temp5678[22]) );
  DFFQXL \temp5678_reg[21]  ( .D(N181), .CK(clk), .Q(temp5678[21]) );
  DFFQXL \temp5678_reg[20]  ( .D(N180), .CK(clk), .Q(temp5678[20]) );
  DFFQXL \temp34_reg[26]  ( .D(N58), .CK(clk), .Q(temp34[26]) );
  DFFQXL \temp34_reg[25]  ( .D(N57), .CK(clk), .Q(temp34[25]) );
  DFFQXL \temp34_reg[24]  ( .D(N56), .CK(clk), .Q(temp34[24]) );
  DFFQXL \temp34_reg[23]  ( .D(N55), .CK(clk), .Q(temp34[23]) );
  DFFQXL \temp34_reg[22]  ( .D(N54), .CK(clk), .Q(temp34[22]) );
  DFFQXL \temp34_reg[21]  ( .D(N53), .CK(clk), .Q(temp34[21]) );
  DFFQXL \temp34_reg[20]  ( .D(N52), .CK(clk), .Q(temp34[20]) );
  DFFQXL \temp78_reg[26]  ( .D(N122), .CK(clk), .Q(temp78[26]) );
  DFFQXL \temp78_reg[25]  ( .D(N121), .CK(clk), .Q(temp78[25]) );
  DFFQXL \temp78_reg[24]  ( .D(N120), .CK(clk), .Q(temp78[24]) );
  DFFQXL \temp78_reg[23]  ( .D(N119), .CK(clk), .Q(temp78[23]) );
  DFFQXL \temp78_reg[22]  ( .D(N118), .CK(clk), .Q(temp78[22]) );
  DFFQXL \temp78_reg[21]  ( .D(N117), .CK(clk), .Q(temp78[21]) );
  DFFQXL \temp78_reg[20]  ( .D(N116), .CK(clk), .Q(temp78[20]) );
  DFFQXL \temp1234_reg[28]  ( .D(N156), .CK(clk), .Q(temp1234[28]) );
  DFFQXL \temp1234_reg[27]  ( .D(N155), .CK(clk), .Q(temp1234[27]) );
  DFFQXL \temp1234_reg[26]  ( .D(N154), .CK(clk), .Q(temp1234[26]) );
  DFFQXL \temp1234_reg[25]  ( .D(N153), .CK(clk), .Q(temp1234[25]) );
  DFFQXL \temp1234_reg[24]  ( .D(N152), .CK(clk), .Q(temp1234[24]) );
  DFFQXL \temp1234_reg[23]  ( .D(N151), .CK(clk), .Q(temp1234[23]) );
  DFFQXL \temp1234_reg[22]  ( .D(N150), .CK(clk), .Q(temp1234[22]) );
  DFFQXL \temp1234_reg[21]  ( .D(N149), .CK(clk), .Q(temp1234[21]) );
  DFFQXL \temp9_2_reg[21]  ( .D(temp9[21]), .CK(clk), .Q(temp9_2[21]) );
  DFFQXL \temp9_2_reg[20]  ( .D(temp9[20]), .CK(clk), .Q(temp9_2[20]) );
  DFFQXL \temp9_2_reg[19]  ( .D(temp9[19]), .CK(clk), .Q(temp9_2[19]) );
  DFFQXL \temp9_2_reg[18]  ( .D(temp9[18]), .CK(clk), .Q(temp9_2[18]) );
  DFFQXL \temp9_2_reg[17]  ( .D(temp9[17]), .CK(clk), .Q(temp9_2[17]) );
  DFFQXL \temp9_2_reg[16]  ( .D(temp9[16]), .CK(clk), .Q(temp9_2[16]) );
  DFFQXL \temp9_2_reg[15]  ( .D(temp9[15]), .CK(clk), .Q(temp9_2[15]) );
  DFFQXL \temp9_2_reg[14]  ( .D(temp9[14]), .CK(clk), .Q(temp9_2[14]) );
  DFFQXL \temp12_reg[19]  ( .D(N19), .CK(clk), .Q(temp12[19]) );
  DFFQXL \temp12_reg[18]  ( .D(N18), .CK(clk), .Q(temp12[18]) );
  DFFQXL \temp12_reg[17]  ( .D(N17), .CK(clk), .Q(temp12[17]) );
  DFFQXL \temp12_reg[16]  ( .D(N16), .CK(clk), .Q(temp12[16]) );
  DFFQXL \temp12_reg[15]  ( .D(N15), .CK(clk), .Q(temp12[15]) );
  DFFQXL \temp12_reg[14]  ( .D(N14), .CK(clk), .Q(temp12[14]) );
  DFFQXL \temp12_reg[13]  ( .D(N13), .CK(clk), .Q(temp12[13]) );
  DFFQXL \temp12_reg[12]  ( .D(N12), .CK(clk), .Q(temp12[12]) );
  DFFQXL \temp56_reg[19]  ( .D(N83), .CK(clk), .Q(temp56[19]) );
  DFFQXL \temp56_reg[18]  ( .D(N82), .CK(clk), .Q(temp56[18]) );
  DFFQXL \temp56_reg[17]  ( .D(N81), .CK(clk), .Q(temp56[17]) );
  DFFQXL \temp56_reg[16]  ( .D(N80), .CK(clk), .Q(temp56[16]) );
  DFFQXL \temp56_reg[15]  ( .D(N79), .CK(clk), .Q(temp56[15]) );
  DFFQXL \temp56_reg[14]  ( .D(N78), .CK(clk), .Q(temp56[14]) );
  DFFQXL \temp56_reg[13]  ( .D(N77), .CK(clk), .Q(temp56[13]) );
  DFFQXL \temp56_reg[12]  ( .D(N76), .CK(clk), .Q(temp56[12]) );
  DFFQXL \temp5678_reg[19]  ( .D(N179), .CK(clk), .Q(temp5678[19]) );
  DFFQXL \temp5678_reg[18]  ( .D(N178), .CK(clk), .Q(temp5678[18]) );
  DFFQXL \temp5678_reg[17]  ( .D(N177), .CK(clk), .Q(temp5678[17]) );
  DFFQXL \temp5678_reg[16]  ( .D(N176), .CK(clk), .Q(temp5678[16]) );
  DFFQXL \temp5678_reg[15]  ( .D(N175), .CK(clk), .Q(temp5678[15]) );
  DFFQXL \temp5678_reg[14]  ( .D(N174), .CK(clk), .Q(temp5678[14]) );
  DFFQXL \temp5678_reg[13]  ( .D(N173), .CK(clk), .Q(temp5678[13]) );
  DFFQXL \temp5678_reg[12]  ( .D(N172), .CK(clk), .Q(temp5678[12]) );
  DFFQXL \temp34_reg[19]  ( .D(N51), .CK(clk), .Q(temp34[19]) );
  DFFQXL \temp34_reg[18]  ( .D(N50), .CK(clk), .Q(temp34[18]) );
  DFFQXL \temp34_reg[17]  ( .D(N49), .CK(clk), .Q(temp34[17]) );
  DFFQXL \temp34_reg[16]  ( .D(N48), .CK(clk), .Q(temp34[16]) );
  DFFQXL \temp34_reg[15]  ( .D(N47), .CK(clk), .Q(temp34[15]) );
  DFFQXL \temp34_reg[14]  ( .D(N46), .CK(clk), .Q(temp34[14]) );
  DFFQXL \temp34_reg[13]  ( .D(N45), .CK(clk), .Q(temp34[13]) );
  DFFQXL \temp34_reg[12]  ( .D(N44), .CK(clk), .Q(temp34[12]) );
  DFFQXL \temp78_reg[19]  ( .D(N115), .CK(clk), .Q(temp78[19]) );
  DFFQXL \temp78_reg[18]  ( .D(N114), .CK(clk), .Q(temp78[18]) );
  DFFQXL \temp78_reg[17]  ( .D(N113), .CK(clk), .Q(temp78[17]) );
  DFFQXL \temp78_reg[16]  ( .D(N112), .CK(clk), .Q(temp78[16]) );
  DFFQXL \temp78_reg[15]  ( .D(N111), .CK(clk), .Q(temp78[15]) );
  DFFQXL \temp78_reg[14]  ( .D(N110), .CK(clk), .Q(temp78[14]) );
  DFFQXL \temp78_reg[13]  ( .D(N109), .CK(clk), .Q(temp78[13]) );
  DFFQXL \temp78_reg[12]  ( .D(N108), .CK(clk), .Q(temp78[12]) );
  DFFQXL \temp1234_reg[20]  ( .D(N148), .CK(clk), .Q(temp1234[20]) );
  DFFQXL \temp1234_reg[19]  ( .D(N147), .CK(clk), .Q(temp1234[19]) );
  DFFQXL \temp1234_reg[18]  ( .D(N146), .CK(clk), .Q(temp1234[18]) );
  DFFQXL \temp1234_reg[17]  ( .D(N145), .CK(clk), .Q(temp1234[17]) );
  DFFQXL \temp1234_reg[16]  ( .D(N144), .CK(clk), .Q(temp1234[16]) );
  DFFQXL \temp1234_reg[15]  ( .D(N143), .CK(clk), .Q(temp1234[15]) );
  DFFQXL \temp1234_reg[14]  ( .D(N142), .CK(clk), .Q(temp1234[14]) );
  DFFQXL \temp9_2_reg[13]  ( .D(temp9[13]), .CK(clk), .Q(temp9_2[13]) );
  DFFQXL \temp9_2_reg[12]  ( .D(temp9[12]), .CK(clk), .Q(temp9_2[12]) );
  DFFQXL \temp9_2_reg[11]  ( .D(temp9[11]), .CK(clk), .Q(temp9_2[11]) );
  DFFQXL \temp9_2_reg[10]  ( .D(temp9[10]), .CK(clk), .Q(temp9_2[10]) );
  DFFQXL \temp9_2_reg[9]  ( .D(temp9[9]), .CK(clk), .Q(temp9_2[9]) );
  DFFQXL \temp9_2_reg[8]  ( .D(temp9[8]), .CK(clk), .Q(temp9_2[8]) );
  DFFQXL \temp9_2_reg[7]  ( .D(temp9[7]), .CK(clk), .Q(temp9_2[7]) );
  DFFQXL \temp12_reg[11]  ( .D(N11), .CK(clk), .Q(temp12[11]) );
  DFFQXL \temp12_reg[10]  ( .D(N10), .CK(clk), .Q(temp12[10]) );
  DFFQXL \temp12_reg[9]  ( .D(N9), .CK(clk), .Q(temp12[9]) );
  DFFQXL \temp12_reg[8]  ( .D(N8), .CK(clk), .Q(temp12[8]) );
  DFFQXL \temp12_reg[7]  ( .D(N7), .CK(clk), .Q(temp12[7]) );
  DFFQXL \temp12_reg[6]  ( .D(N6), .CK(clk), .Q(temp12[6]) );
  DFFQXL \temp12_reg[5]  ( .D(N5), .CK(clk), .Q(temp12[5]) );
  DFFQXL \temp56_reg[11]  ( .D(N75), .CK(clk), .Q(temp56[11]) );
  DFFQXL \temp56_reg[10]  ( .D(N74), .CK(clk), .Q(temp56[10]) );
  DFFQXL \temp56_reg[9]  ( .D(N73), .CK(clk), .Q(temp56[9]) );
  DFFQXL \temp56_reg[8]  ( .D(N72), .CK(clk), .Q(temp56[8]) );
  DFFQXL \temp56_reg[7]  ( .D(N71), .CK(clk), .Q(temp56[7]) );
  DFFQXL \temp56_reg[6]  ( .D(N70), .CK(clk), .Q(temp56[6]) );
  DFFQXL \temp56_reg[5]  ( .D(N69), .CK(clk), .Q(temp56[5]) );
  DFFQXL \temp5678_reg[11]  ( .D(N171), .CK(clk), .Q(temp5678[11]) );
  DFFQXL \temp5678_reg[10]  ( .D(N170), .CK(clk), .Q(temp5678[10]) );
  DFFQXL \temp5678_reg[9]  ( .D(N169), .CK(clk), .Q(temp5678[9]) );
  DFFQXL \temp5678_reg[8]  ( .D(N168), .CK(clk), .Q(temp5678[8]) );
  DFFQXL \temp5678_reg[7]  ( .D(N167), .CK(clk), .Q(temp5678[7]) );
  DFFQXL \temp5678_reg[6]  ( .D(N166), .CK(clk), .Q(temp5678[6]) );
  DFFQXL \temp5678_reg[5]  ( .D(N165), .CK(clk), .Q(temp5678[5]) );
  DFFQXL \temp34_reg[11]  ( .D(N43), .CK(clk), .Q(temp34[11]) );
  DFFQXL \temp34_reg[10]  ( .D(N42), .CK(clk), .Q(temp34[10]) );
  DFFQXL \temp34_reg[9]  ( .D(N41), .CK(clk), .Q(temp34[9]) );
  DFFQXL \temp34_reg[8]  ( .D(N40), .CK(clk), .Q(temp34[8]) );
  DFFQXL \temp34_reg[7]  ( .D(N39), .CK(clk), .Q(temp34[7]) );
  DFFQXL \temp34_reg[6]  ( .D(N38), .CK(clk), .Q(temp34[6]) );
  DFFQXL \temp34_reg[5]  ( .D(N37), .CK(clk), .Q(temp34[5]) );
  DFFQXL \temp78_reg[11]  ( .D(N107), .CK(clk), .Q(temp78[11]) );
  DFFQXL \temp78_reg[10]  ( .D(N106), .CK(clk), .Q(temp78[10]) );
  DFFQXL \temp78_reg[9]  ( .D(N105), .CK(clk), .Q(temp78[9]) );
  DFFQXL \temp78_reg[8]  ( .D(N104), .CK(clk), .Q(temp78[8]) );
  DFFQXL \temp78_reg[7]  ( .D(N103), .CK(clk), .Q(temp78[7]) );
  DFFQXL \temp78_reg[6]  ( .D(N102), .CK(clk), .Q(temp78[6]) );
  DFFQXL \temp78_reg[5]  ( .D(N101), .CK(clk), .Q(temp78[5]) );
  DFFQXL \temp1234_reg[13]  ( .D(N141), .CK(clk), .Q(temp1234[13]) );
  DFFQXL \temp1234_reg[12]  ( .D(N140), .CK(clk), .Q(temp1234[12]) );
  DFFQXL \temp1234_reg[11]  ( .D(N139), .CK(clk), .Q(temp1234[11]) );
  DFFQXL \temp1234_reg[10]  ( .D(N138), .CK(clk), .Q(temp1234[10]) );
  DFFQXL \temp1234_reg[9]  ( .D(N137), .CK(clk), .Q(temp1234[9]) );
  DFFQXL \temp1234_reg[8]  ( .D(N136), .CK(clk), .Q(temp1234[8]) );
  DFFQXL \temp1234_reg[7]  ( .D(N135), .CK(clk), .Q(temp1234[7]) );
  DFFQXL \temp1234_reg[6]  ( .D(N134), .CK(clk), .Q(temp1234[6]) );
  DFFQXL \temp9_2_reg[6]  ( .D(temp9[6]), .CK(clk), .Q(temp9_2[6]) );
  DFFQXL \temp9_2_reg[5]  ( .D(temp9[5]), .CK(clk), .Q(temp9_2[5]) );
  DFFQXL \temp9_2_reg[4]  ( .D(temp9[4]), .CK(clk), .Q(temp9_2[4]) );
  DFFQXL \temp9_2_reg[3]  ( .D(temp9[3]), .CK(clk), .Q(temp9_2[3]) );
  DFFQXL \temp9_2_reg[2]  ( .D(temp9[2]), .CK(clk), .Q(temp9_2[2]) );
  DFFQXL \temp9_2_reg[1]  ( .D(temp9[1]), .CK(clk), .Q(temp9_2[1]) );
  DFFQXL \temp12_reg[4]  ( .D(N4), .CK(clk), .Q(temp12[4]) );
  DFFQXL \temp12_reg[3]  ( .D(N3), .CK(clk), .Q(temp12[3]) );
  DFFQXL \temp12_reg[2]  ( .D(N2), .CK(clk), .Q(temp12[2]) );
  DFFQXL \temp12_reg[1]  ( .D(N1), .CK(clk), .Q(temp12[1]) );
  DFFQXL \temp56_reg[4]  ( .D(N68), .CK(clk), .Q(temp56[4]) );
  DFFQXL \temp56_reg[3]  ( .D(N67), .CK(clk), .Q(temp56[3]) );
  DFFQXL \temp56_reg[2]  ( .D(N66), .CK(clk), .Q(temp56[2]) );
  DFFQXL \temp56_reg[1]  ( .D(N65), .CK(clk), .Q(temp56[1]) );
  DFFQXL \temp5678_reg[4]  ( .D(N164), .CK(clk), .Q(temp5678[4]) );
  DFFQXL \temp5678_reg[3]  ( .D(N163), .CK(clk), .Q(temp5678[3]) );
  DFFQXL \temp5678_reg[2]  ( .D(N162), .CK(clk), .Q(temp5678[2]) );
  DFFQXL \temp5678_reg[1]  ( .D(N161), .CK(clk), .Q(temp5678[1]) );
  DFFQXL \temp34_reg[4]  ( .D(N36), .CK(clk), .Q(temp34[4]) );
  DFFQXL \temp34_reg[3]  ( .D(N35), .CK(clk), .Q(temp34[3]) );
  DFFQXL \temp34_reg[2]  ( .D(N34), .CK(clk), .Q(temp34[2]) );
  DFFQXL \temp34_reg[1]  ( .D(N33), .CK(clk), .Q(temp34[1]) );
  DFFQXL \temp78_reg[4]  ( .D(N100), .CK(clk), .Q(temp78[4]) );
  DFFQXL \temp78_reg[3]  ( .D(N99), .CK(clk), .Q(temp78[3]) );
  DFFQXL \temp78_reg[2]  ( .D(N98), .CK(clk), .Q(temp78[2]) );
  DFFQXL \temp78_reg[1]  ( .D(N97), .CK(clk), .Q(temp78[1]) );
  DFFQXL \temp1234_reg[5]  ( .D(N133), .CK(clk), .Q(temp1234[5]) );
  DFFQXL \temp1234_reg[4]  ( .D(N132), .CK(clk), .Q(temp1234[4]) );
  DFFQXL \temp1234_reg[3]  ( .D(N131), .CK(clk), .Q(temp1234[3]) );
  DFFQXL \temp1234_reg[2]  ( .D(N130), .CK(clk), .Q(temp1234[2]) );
  DFFQXL \temp1234_reg[1]  ( .D(N129), .CK(clk), .Q(temp1234[1]) );
  DFFQXL \total_reg[31]  ( .D(N255), .CK(clk), .Q(total[31]) );
  DFFQXL \total_reg[30]  ( .D(N254), .CK(clk), .Q(total[30]) );
  DFFQXL \total_reg[29]  ( .D(N253), .CK(clk), .Q(total[29]) );
  DFFQXL \total_reg[28]  ( .D(N252), .CK(clk), .Q(total[28]) );
  DFFQXL \total_reg[27]  ( .D(N251), .CK(clk), .Q(total[27]) );
  DFFQXL \total_reg[26]  ( .D(N250), .CK(clk), .Q(total[26]) );
  DFFQXL \total_reg[25]  ( .D(N249), .CK(clk), .Q(total[25]) );
  DFFQXL \total_reg[24]  ( .D(N248), .CK(clk), .Q(total[24]) );
  DFFQXL \total_reg[23]  ( .D(N247), .CK(clk), .Q(total[23]) );
  DFFQXL \total_reg[22]  ( .D(N246), .CK(clk), .Q(total[22]) );
  DFFQXL \total_reg[21]  ( .D(N245), .CK(clk), .Q(total[21]) );
  DFFQXL \total_reg[20]  ( .D(N244), .CK(clk), .Q(total[20]) );
  DFFQXL \total_reg[19]  ( .D(N243), .CK(clk), .Q(total[19]) );
  DFFQXL \total_reg[18]  ( .D(N242), .CK(clk), .Q(total[18]) );
  DFFQXL \total_reg[17]  ( .D(N241), .CK(clk), .Q(total[17]) );
  DFFQXL \total_reg[16]  ( .D(N240), .CK(clk), .Q(total[16]) );
  DFFQXL \total_reg[15]  ( .D(N239), .CK(clk), .Q(total[15]) );
  DFFQXL \total_reg[14]  ( .D(N238), .CK(clk), .Q(total[14]) );
  DFFQXL \total_reg[13]  ( .D(N237), .CK(clk), .Q(total[13]) );
  DFFQXL \total_reg[12]  ( .D(N236), .CK(clk), .Q(total[12]) );
  DFFQXL \total_reg[11]  ( .D(N235), .CK(clk), .Q(total[11]) );
  DFFQXL \total_reg[10]  ( .D(N234), .CK(clk), .Q(total[10]) );
  DFFQXL \total_reg[9]  ( .D(N233), .CK(clk), .Q(total[9]) );
  DFFQXL \total_reg[8]  ( .D(N232), .CK(clk), .Q(total[8]) );
  DFFQXL \total_reg[7]  ( .D(N231), .CK(clk), .Q(total[7]) );
  DFFQXL \total_reg[6]  ( .D(N230), .CK(clk), .Q(total[6]) );
  DFFQXL \total_reg[5]  ( .D(N229), .CK(clk), .Q(total[5]) );
  DFFQXL \total_reg[4]  ( .D(N228), .CK(clk), .Q(total[4]) );
  DFFQXL \total_reg[3]  ( .D(N227), .CK(clk), .Q(total[3]) );
  DFFQXL \total_reg[2]  ( .D(N226), .CK(clk), .Q(total[2]) );
  DFFQXL \total_reg[1]  ( .D(N225), .CK(clk), .Q(total[1]) );
  DFFQXL \total_reg[0]  ( .D(N224), .CK(clk), .Q(total[0]) );
  DFFQXL \temp34_reg[0]  ( .D(N32), .CK(clk), .Q(temp34[0]) );
  DFFQXL \temp78_reg[0]  ( .D(N96), .CK(clk), .Q(temp78[0]) );
  DFFQXL \temp1234_reg[0]  ( .D(N128), .CK(clk), .Q(temp1234[0]) );
  DFFQXL \temp12_reg[0]  ( .D(N0), .CK(clk), .Q(temp12[0]) );
  DFFQXL \temp56_reg[0]  ( .D(N64), .CK(clk), .Q(temp56[0]) );
  DFFQXL \temp5678_reg[0]  ( .D(N160), .CK(clk), .Q(temp5678[0]) );
  DFFQXL \temp9_2_reg[0]  ( .D(temp9[0]), .CK(clk), .Q(temp9_2[0]) );
  DFFQXL \temp9_reg[31]  ( .D(in9[31]), .CK(clk), .Q(temp9[31]) );
  DFFQXL \temp9_reg[30]  ( .D(in9[30]), .CK(clk), .Q(temp9[30]) );
  DFFQXL \temp9_reg[29]  ( .D(in9[29]), .CK(clk), .Q(temp9[29]) );
  DFFQXL \temp9_reg[28]  ( .D(in9[28]), .CK(clk), .Q(temp9[28]) );
  DFFQXL \temp9_reg[27]  ( .D(in9[27]), .CK(clk), .Q(temp9[27]) );
  DFFQXL \temp9_reg[26]  ( .D(in9[26]), .CK(clk), .Q(temp9[26]) );
  DFFQXL \temp9_reg[25]  ( .D(in9[25]), .CK(clk), .Q(temp9[25]) );
  DFFQXL \temp9_reg[24]  ( .D(in9[24]), .CK(clk), .Q(temp9[24]) );
  DFFQXL \temp9_reg[23]  ( .D(in9[23]), .CK(clk), .Q(temp9[23]) );
  DFFQXL \temp9_reg[22]  ( .D(in9[22]), .CK(clk), .Q(temp9[22]) );
  DFFQXL \temp9_reg[21]  ( .D(in9[21]), .CK(clk), .Q(temp9[21]) );
  DFFQXL \temp9_reg[20]  ( .D(in9[20]), .CK(clk), .Q(temp9[20]) );
  DFFQXL \temp9_reg[19]  ( .D(in9[19]), .CK(clk), .Q(temp9[19]) );
  DFFQXL \temp9_reg[18]  ( .D(in9[18]), .CK(clk), .Q(temp9[18]) );
  DFFQXL \temp9_reg[17]  ( .D(in9[17]), .CK(clk), .Q(temp9[17]) );
  DFFQXL \temp9_reg[16]  ( .D(in9[16]), .CK(clk), .Q(temp9[16]) );
  DFFQXL \temp9_reg[15]  ( .D(in9[15]), .CK(clk), .Q(temp9[15]) );
  DFFQXL \temp9_reg[14]  ( .D(in9[14]), .CK(clk), .Q(temp9[14]) );
  DFFQXL \temp9_reg[13]  ( .D(in9[13]), .CK(clk), .Q(temp9[13]) );
  DFFQXL \temp9_reg[12]  ( .D(in9[12]), .CK(clk), .Q(temp9[12]) );
  DFFQXL \temp9_reg[11]  ( .D(in9[11]), .CK(clk), .Q(temp9[11]) );
  DFFQXL \temp9_reg[10]  ( .D(in9[10]), .CK(clk), .Q(temp9[10]) );
  DFFQXL \temp9_reg[9]  ( .D(in9[9]), .CK(clk), .Q(temp9[9]) );
  DFFQXL \temp9_reg[8]  ( .D(in9[8]), .CK(clk), .Q(temp9[8]) );
  DFFQXL \temp9_reg[7]  ( .D(in9[7]), .CK(clk), .Q(temp9[7]) );
  DFFQXL \temp9_reg[6]  ( .D(in9[6]), .CK(clk), .Q(temp9[6]) );
  DFFQXL \temp9_reg[5]  ( .D(in9[5]), .CK(clk), .Q(temp9[5]) );
  DFFQXL \temp9_reg[4]  ( .D(in9[4]), .CK(clk), .Q(temp9[4]) );
  DFFQXL \temp9_reg[3]  ( .D(in9[3]), .CK(clk), .Q(temp9[3]) );
  DFFQXL \temp9_reg[2]  ( .D(in9[2]), .CK(clk), .Q(temp9[2]) );
  DFFQXL \temp9_reg[1]  ( .D(in9[1]), .CK(clk), .Q(temp9[1]) );
  DFFQXL \temp9_reg[0]  ( .D(in9[0]), .CK(clk), .Q(temp9[0]) );
endmodule


module Adder_tree_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_2 ( in1, in2, in3, in4, in5, in6, in7, in8, in9, total, clk
 );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  input [31:0] in5;
  input [31:0] in6;
  input [31:0] in7;
  input [31:0] in8;
  input [31:0] in9;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N223, N222, N221, N220, N219, N218, N217, N216,
         N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205,
         N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194,
         N193, N192;
  wire   [31:0] temp9;
  wire   [31:0] temp12;
  wire   [31:0] temp34;
  wire   [31:0] temp56;
  wire   [31:0] temp78;
  wire   [31:0] temp1234;
  wire   [31:0] temp5678;
  wire   [31:0] temp9_2;

  Adder_tree_2_DW01_add_0 add_29 ( .A(temp56), .B(temp78), .CI(1'b0), .SUM({
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160}) );
  Adder_tree_2_DW01_add_1 add_28 ( .A(temp12), .B(temp34), .CI(1'b0), .SUM({
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, 
        N135, N134, N133, N132, N131, N130, N129, N128}) );
  Adder_tree_2_DW01_add_2 add_25 ( .A(in7), .B(in8), .CI(1'b0), .SUM({N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96}) );
  Adder_tree_2_DW01_add_3 add_24 ( .A(in5), .B(in6), .CI(1'b0), .SUM({N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64}) );
  Adder_tree_2_DW01_add_4 add_23 ( .A(in3), .B(in4), .CI(1'b0), .SUM({N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32}) );
  Adder_tree_2_DW01_add_5 add_22 ( .A(in1), .B(in2), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Adder_tree_2_DW01_add_7 add_1_root_add_0_root_add_32_2 ( .A(temp9_2), .B(
        temp1234), .CI(1'b0), .SUM({N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 
        N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, 
        N192}) );
  Adder_tree_2_DW01_add_6 add_0_root_add_0_root_add_32_2 ( .A(temp5678), .B({
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192}), .CI(1'b0), .SUM({
        N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, 
        N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, 
        N231, N230, N229, N228, N227, N226, N225, N224}) );
  DFFQXL \temp9_2_reg[31]  ( .D(temp9[31]), .CK(clk), .Q(temp9_2[31]) );
  DFFQXL \temp9_2_reg[30]  ( .D(temp9[30]), .CK(clk), .Q(temp9_2[30]) );
  DFFQXL \temp9_2_reg[29]  ( .D(temp9[29]), .CK(clk), .Q(temp9_2[29]) );
  DFFQXL \temp12_reg[31]  ( .D(N31), .CK(clk), .Q(temp12[31]) );
  DFFQXL \temp12_reg[30]  ( .D(N30), .CK(clk), .Q(temp12[30]) );
  DFFQXL \temp12_reg[29]  ( .D(N29), .CK(clk), .Q(temp12[29]) );
  DFFQXL \temp12_reg[28]  ( .D(N28), .CK(clk), .Q(temp12[28]) );
  DFFQXL \temp12_reg[27]  ( .D(N27), .CK(clk), .Q(temp12[27]) );
  DFFQXL \temp56_reg[31]  ( .D(N95), .CK(clk), .Q(temp56[31]) );
  DFFQXL \temp56_reg[30]  ( .D(N94), .CK(clk), .Q(temp56[30]) );
  DFFQXL \temp56_reg[29]  ( .D(N93), .CK(clk), .Q(temp56[29]) );
  DFFQXL \temp56_reg[28]  ( .D(N92), .CK(clk), .Q(temp56[28]) );
  DFFQXL \temp56_reg[27]  ( .D(N91), .CK(clk), .Q(temp56[27]) );
  DFFQXL \temp5678_reg[31]  ( .D(N191), .CK(clk), .Q(temp5678[31]) );
  DFFQXL \temp5678_reg[30]  ( .D(N190), .CK(clk), .Q(temp5678[30]) );
  DFFQXL \temp5678_reg[29]  ( .D(N189), .CK(clk), .Q(temp5678[29]) );
  DFFQXL \temp5678_reg[28]  ( .D(N188), .CK(clk), .Q(temp5678[28]) );
  DFFQXL \temp5678_reg[27]  ( .D(N187), .CK(clk), .Q(temp5678[27]) );
  DFFQXL \temp34_reg[31]  ( .D(N63), .CK(clk), .Q(temp34[31]) );
  DFFQXL \temp34_reg[30]  ( .D(N62), .CK(clk), .Q(temp34[30]) );
  DFFQXL \temp34_reg[29]  ( .D(N61), .CK(clk), .Q(temp34[29]) );
  DFFQXL \temp34_reg[28]  ( .D(N60), .CK(clk), .Q(temp34[28]) );
  DFFQXL \temp34_reg[27]  ( .D(N59), .CK(clk), .Q(temp34[27]) );
  DFFQXL \temp78_reg[31]  ( .D(N127), .CK(clk), .Q(temp78[31]) );
  DFFQXL \temp78_reg[30]  ( .D(N126), .CK(clk), .Q(temp78[30]) );
  DFFQXL \temp78_reg[29]  ( .D(N125), .CK(clk), .Q(temp78[29]) );
  DFFQXL \temp78_reg[28]  ( .D(N124), .CK(clk), .Q(temp78[28]) );
  DFFQXL \temp78_reg[27]  ( .D(N123), .CK(clk), .Q(temp78[27]) );
  DFFQXL \temp1234_reg[31]  ( .D(N159), .CK(clk), .Q(temp1234[31]) );
  DFFQXL \temp1234_reg[30]  ( .D(N158), .CK(clk), .Q(temp1234[30]) );
  DFFQXL \temp1234_reg[29]  ( .D(N157), .CK(clk), .Q(temp1234[29]) );
  DFFQXL \temp9_2_reg[28]  ( .D(temp9[28]), .CK(clk), .Q(temp9_2[28]) );
  DFFQXL \temp9_2_reg[27]  ( .D(temp9[27]), .CK(clk), .Q(temp9_2[27]) );
  DFFQXL \temp9_2_reg[26]  ( .D(temp9[26]), .CK(clk), .Q(temp9_2[26]) );
  DFFQXL \temp9_2_reg[25]  ( .D(temp9[25]), .CK(clk), .Q(temp9_2[25]) );
  DFFQXL \temp9_2_reg[24]  ( .D(temp9[24]), .CK(clk), .Q(temp9_2[24]) );
  DFFQXL \temp9_2_reg[23]  ( .D(temp9[23]), .CK(clk), .Q(temp9_2[23]) );
  DFFQXL \temp9_2_reg[22]  ( .D(temp9[22]), .CK(clk), .Q(temp9_2[22]) );
  DFFQXL \temp12_reg[26]  ( .D(N26), .CK(clk), .Q(temp12[26]) );
  DFFQXL \temp12_reg[25]  ( .D(N25), .CK(clk), .Q(temp12[25]) );
  DFFQXL \temp12_reg[24]  ( .D(N24), .CK(clk), .Q(temp12[24]) );
  DFFQXL \temp12_reg[23]  ( .D(N23), .CK(clk), .Q(temp12[23]) );
  DFFQXL \temp12_reg[22]  ( .D(N22), .CK(clk), .Q(temp12[22]) );
  DFFQXL \temp12_reg[21]  ( .D(N21), .CK(clk), .Q(temp12[21]) );
  DFFQXL \temp12_reg[20]  ( .D(N20), .CK(clk), .Q(temp12[20]) );
  DFFQXL \temp56_reg[26]  ( .D(N90), .CK(clk), .Q(temp56[26]) );
  DFFQXL \temp56_reg[25]  ( .D(N89), .CK(clk), .Q(temp56[25]) );
  DFFQXL \temp56_reg[24]  ( .D(N88), .CK(clk), .Q(temp56[24]) );
  DFFQXL \temp56_reg[23]  ( .D(N87), .CK(clk), .Q(temp56[23]) );
  DFFQXL \temp56_reg[22]  ( .D(N86), .CK(clk), .Q(temp56[22]) );
  DFFQXL \temp56_reg[21]  ( .D(N85), .CK(clk), .Q(temp56[21]) );
  DFFQXL \temp56_reg[20]  ( .D(N84), .CK(clk), .Q(temp56[20]) );
  DFFQXL \temp5678_reg[26]  ( .D(N186), .CK(clk), .Q(temp5678[26]) );
  DFFQXL \temp5678_reg[25]  ( .D(N185), .CK(clk), .Q(temp5678[25]) );
  DFFQXL \temp5678_reg[24]  ( .D(N184), .CK(clk), .Q(temp5678[24]) );
  DFFQXL \temp5678_reg[23]  ( .D(N183), .CK(clk), .Q(temp5678[23]) );
  DFFQXL \temp5678_reg[22]  ( .D(N182), .CK(clk), .Q(temp5678[22]) );
  DFFQXL \temp5678_reg[21]  ( .D(N181), .CK(clk), .Q(temp5678[21]) );
  DFFQXL \temp5678_reg[20]  ( .D(N180), .CK(clk), .Q(temp5678[20]) );
  DFFQXL \temp34_reg[26]  ( .D(N58), .CK(clk), .Q(temp34[26]) );
  DFFQXL \temp34_reg[25]  ( .D(N57), .CK(clk), .Q(temp34[25]) );
  DFFQXL \temp34_reg[24]  ( .D(N56), .CK(clk), .Q(temp34[24]) );
  DFFQXL \temp34_reg[23]  ( .D(N55), .CK(clk), .Q(temp34[23]) );
  DFFQXL \temp34_reg[22]  ( .D(N54), .CK(clk), .Q(temp34[22]) );
  DFFQXL \temp34_reg[21]  ( .D(N53), .CK(clk), .Q(temp34[21]) );
  DFFQXL \temp34_reg[20]  ( .D(N52), .CK(clk), .Q(temp34[20]) );
  DFFQXL \temp78_reg[26]  ( .D(N122), .CK(clk), .Q(temp78[26]) );
  DFFQXL \temp78_reg[25]  ( .D(N121), .CK(clk), .Q(temp78[25]) );
  DFFQXL \temp78_reg[24]  ( .D(N120), .CK(clk), .Q(temp78[24]) );
  DFFQXL \temp78_reg[23]  ( .D(N119), .CK(clk), .Q(temp78[23]) );
  DFFQXL \temp78_reg[22]  ( .D(N118), .CK(clk), .Q(temp78[22]) );
  DFFQXL \temp78_reg[21]  ( .D(N117), .CK(clk), .Q(temp78[21]) );
  DFFQXL \temp78_reg[20]  ( .D(N116), .CK(clk), .Q(temp78[20]) );
  DFFQXL \temp1234_reg[28]  ( .D(N156), .CK(clk), .Q(temp1234[28]) );
  DFFQXL \temp1234_reg[27]  ( .D(N155), .CK(clk), .Q(temp1234[27]) );
  DFFQXL \temp1234_reg[26]  ( .D(N154), .CK(clk), .Q(temp1234[26]) );
  DFFQXL \temp1234_reg[25]  ( .D(N153), .CK(clk), .Q(temp1234[25]) );
  DFFQXL \temp1234_reg[24]  ( .D(N152), .CK(clk), .Q(temp1234[24]) );
  DFFQXL \temp1234_reg[23]  ( .D(N151), .CK(clk), .Q(temp1234[23]) );
  DFFQXL \temp1234_reg[22]  ( .D(N150), .CK(clk), .Q(temp1234[22]) );
  DFFQXL \temp1234_reg[21]  ( .D(N149), .CK(clk), .Q(temp1234[21]) );
  DFFQXL \temp9_2_reg[21]  ( .D(temp9[21]), .CK(clk), .Q(temp9_2[21]) );
  DFFQXL \temp9_2_reg[20]  ( .D(temp9[20]), .CK(clk), .Q(temp9_2[20]) );
  DFFQXL \temp9_2_reg[19]  ( .D(temp9[19]), .CK(clk), .Q(temp9_2[19]) );
  DFFQXL \temp9_2_reg[18]  ( .D(temp9[18]), .CK(clk), .Q(temp9_2[18]) );
  DFFQXL \temp9_2_reg[17]  ( .D(temp9[17]), .CK(clk), .Q(temp9_2[17]) );
  DFFQXL \temp9_2_reg[16]  ( .D(temp9[16]), .CK(clk), .Q(temp9_2[16]) );
  DFFQXL \temp9_2_reg[15]  ( .D(temp9[15]), .CK(clk), .Q(temp9_2[15]) );
  DFFQXL \temp9_2_reg[14]  ( .D(temp9[14]), .CK(clk), .Q(temp9_2[14]) );
  DFFQXL \temp12_reg[19]  ( .D(N19), .CK(clk), .Q(temp12[19]) );
  DFFQXL \temp12_reg[18]  ( .D(N18), .CK(clk), .Q(temp12[18]) );
  DFFQXL \temp12_reg[17]  ( .D(N17), .CK(clk), .Q(temp12[17]) );
  DFFQXL \temp12_reg[16]  ( .D(N16), .CK(clk), .Q(temp12[16]) );
  DFFQXL \temp12_reg[15]  ( .D(N15), .CK(clk), .Q(temp12[15]) );
  DFFQXL \temp12_reg[14]  ( .D(N14), .CK(clk), .Q(temp12[14]) );
  DFFQXL \temp12_reg[13]  ( .D(N13), .CK(clk), .Q(temp12[13]) );
  DFFQXL \temp12_reg[12]  ( .D(N12), .CK(clk), .Q(temp12[12]) );
  DFFQXL \temp56_reg[19]  ( .D(N83), .CK(clk), .Q(temp56[19]) );
  DFFQXL \temp56_reg[18]  ( .D(N82), .CK(clk), .Q(temp56[18]) );
  DFFQXL \temp56_reg[17]  ( .D(N81), .CK(clk), .Q(temp56[17]) );
  DFFQXL \temp56_reg[16]  ( .D(N80), .CK(clk), .Q(temp56[16]) );
  DFFQXL \temp56_reg[15]  ( .D(N79), .CK(clk), .Q(temp56[15]) );
  DFFQXL \temp56_reg[14]  ( .D(N78), .CK(clk), .Q(temp56[14]) );
  DFFQXL \temp56_reg[13]  ( .D(N77), .CK(clk), .Q(temp56[13]) );
  DFFQXL \temp56_reg[12]  ( .D(N76), .CK(clk), .Q(temp56[12]) );
  DFFQXL \temp5678_reg[19]  ( .D(N179), .CK(clk), .Q(temp5678[19]) );
  DFFQXL \temp5678_reg[18]  ( .D(N178), .CK(clk), .Q(temp5678[18]) );
  DFFQXL \temp5678_reg[17]  ( .D(N177), .CK(clk), .Q(temp5678[17]) );
  DFFQXL \temp5678_reg[16]  ( .D(N176), .CK(clk), .Q(temp5678[16]) );
  DFFQXL \temp5678_reg[15]  ( .D(N175), .CK(clk), .Q(temp5678[15]) );
  DFFQXL \temp5678_reg[14]  ( .D(N174), .CK(clk), .Q(temp5678[14]) );
  DFFQXL \temp5678_reg[13]  ( .D(N173), .CK(clk), .Q(temp5678[13]) );
  DFFQXL \temp5678_reg[12]  ( .D(N172), .CK(clk), .Q(temp5678[12]) );
  DFFQXL \temp34_reg[19]  ( .D(N51), .CK(clk), .Q(temp34[19]) );
  DFFQXL \temp34_reg[18]  ( .D(N50), .CK(clk), .Q(temp34[18]) );
  DFFQXL \temp34_reg[17]  ( .D(N49), .CK(clk), .Q(temp34[17]) );
  DFFQXL \temp34_reg[16]  ( .D(N48), .CK(clk), .Q(temp34[16]) );
  DFFQXL \temp34_reg[15]  ( .D(N47), .CK(clk), .Q(temp34[15]) );
  DFFQXL \temp34_reg[14]  ( .D(N46), .CK(clk), .Q(temp34[14]) );
  DFFQXL \temp34_reg[13]  ( .D(N45), .CK(clk), .Q(temp34[13]) );
  DFFQXL \temp34_reg[12]  ( .D(N44), .CK(clk), .Q(temp34[12]) );
  DFFQXL \temp78_reg[19]  ( .D(N115), .CK(clk), .Q(temp78[19]) );
  DFFQXL \temp78_reg[18]  ( .D(N114), .CK(clk), .Q(temp78[18]) );
  DFFQXL \temp78_reg[17]  ( .D(N113), .CK(clk), .Q(temp78[17]) );
  DFFQXL \temp78_reg[16]  ( .D(N112), .CK(clk), .Q(temp78[16]) );
  DFFQXL \temp78_reg[15]  ( .D(N111), .CK(clk), .Q(temp78[15]) );
  DFFQXL \temp78_reg[14]  ( .D(N110), .CK(clk), .Q(temp78[14]) );
  DFFQXL \temp78_reg[13]  ( .D(N109), .CK(clk), .Q(temp78[13]) );
  DFFQXL \temp78_reg[12]  ( .D(N108), .CK(clk), .Q(temp78[12]) );
  DFFQXL \temp1234_reg[20]  ( .D(N148), .CK(clk), .Q(temp1234[20]) );
  DFFQXL \temp1234_reg[19]  ( .D(N147), .CK(clk), .Q(temp1234[19]) );
  DFFQXL \temp1234_reg[18]  ( .D(N146), .CK(clk), .Q(temp1234[18]) );
  DFFQXL \temp1234_reg[17]  ( .D(N145), .CK(clk), .Q(temp1234[17]) );
  DFFQXL \temp1234_reg[16]  ( .D(N144), .CK(clk), .Q(temp1234[16]) );
  DFFQXL \temp1234_reg[15]  ( .D(N143), .CK(clk), .Q(temp1234[15]) );
  DFFQXL \temp1234_reg[14]  ( .D(N142), .CK(clk), .Q(temp1234[14]) );
  DFFQXL \temp9_2_reg[13]  ( .D(temp9[13]), .CK(clk), .Q(temp9_2[13]) );
  DFFQXL \temp9_2_reg[12]  ( .D(temp9[12]), .CK(clk), .Q(temp9_2[12]) );
  DFFQXL \temp9_2_reg[11]  ( .D(temp9[11]), .CK(clk), .Q(temp9_2[11]) );
  DFFQXL \temp9_2_reg[10]  ( .D(temp9[10]), .CK(clk), .Q(temp9_2[10]) );
  DFFQXL \temp9_2_reg[9]  ( .D(temp9[9]), .CK(clk), .Q(temp9_2[9]) );
  DFFQXL \temp9_2_reg[8]  ( .D(temp9[8]), .CK(clk), .Q(temp9_2[8]) );
  DFFQXL \temp9_2_reg[7]  ( .D(temp9[7]), .CK(clk), .Q(temp9_2[7]) );
  DFFQXL \temp12_reg[11]  ( .D(N11), .CK(clk), .Q(temp12[11]) );
  DFFQXL \temp12_reg[10]  ( .D(N10), .CK(clk), .Q(temp12[10]) );
  DFFQXL \temp12_reg[9]  ( .D(N9), .CK(clk), .Q(temp12[9]) );
  DFFQXL \temp12_reg[8]  ( .D(N8), .CK(clk), .Q(temp12[8]) );
  DFFQXL \temp12_reg[7]  ( .D(N7), .CK(clk), .Q(temp12[7]) );
  DFFQXL \temp12_reg[6]  ( .D(N6), .CK(clk), .Q(temp12[6]) );
  DFFQXL \temp12_reg[5]  ( .D(N5), .CK(clk), .Q(temp12[5]) );
  DFFQXL \temp56_reg[11]  ( .D(N75), .CK(clk), .Q(temp56[11]) );
  DFFQXL \temp56_reg[10]  ( .D(N74), .CK(clk), .Q(temp56[10]) );
  DFFQXL \temp56_reg[9]  ( .D(N73), .CK(clk), .Q(temp56[9]) );
  DFFQXL \temp56_reg[8]  ( .D(N72), .CK(clk), .Q(temp56[8]) );
  DFFQXL \temp56_reg[7]  ( .D(N71), .CK(clk), .Q(temp56[7]) );
  DFFQXL \temp56_reg[6]  ( .D(N70), .CK(clk), .Q(temp56[6]) );
  DFFQXL \temp56_reg[5]  ( .D(N69), .CK(clk), .Q(temp56[5]) );
  DFFQXL \temp5678_reg[11]  ( .D(N171), .CK(clk), .Q(temp5678[11]) );
  DFFQXL \temp5678_reg[10]  ( .D(N170), .CK(clk), .Q(temp5678[10]) );
  DFFQXL \temp5678_reg[9]  ( .D(N169), .CK(clk), .Q(temp5678[9]) );
  DFFQXL \temp5678_reg[8]  ( .D(N168), .CK(clk), .Q(temp5678[8]) );
  DFFQXL \temp5678_reg[7]  ( .D(N167), .CK(clk), .Q(temp5678[7]) );
  DFFQXL \temp5678_reg[6]  ( .D(N166), .CK(clk), .Q(temp5678[6]) );
  DFFQXL \temp5678_reg[5]  ( .D(N165), .CK(clk), .Q(temp5678[5]) );
  DFFQXL \temp34_reg[11]  ( .D(N43), .CK(clk), .Q(temp34[11]) );
  DFFQXL \temp34_reg[10]  ( .D(N42), .CK(clk), .Q(temp34[10]) );
  DFFQXL \temp34_reg[9]  ( .D(N41), .CK(clk), .Q(temp34[9]) );
  DFFQXL \temp34_reg[8]  ( .D(N40), .CK(clk), .Q(temp34[8]) );
  DFFQXL \temp34_reg[7]  ( .D(N39), .CK(clk), .Q(temp34[7]) );
  DFFQXL \temp34_reg[6]  ( .D(N38), .CK(clk), .Q(temp34[6]) );
  DFFQXL \temp34_reg[5]  ( .D(N37), .CK(clk), .Q(temp34[5]) );
  DFFQXL \temp78_reg[11]  ( .D(N107), .CK(clk), .Q(temp78[11]) );
  DFFQXL \temp78_reg[10]  ( .D(N106), .CK(clk), .Q(temp78[10]) );
  DFFQXL \temp78_reg[9]  ( .D(N105), .CK(clk), .Q(temp78[9]) );
  DFFQXL \temp78_reg[8]  ( .D(N104), .CK(clk), .Q(temp78[8]) );
  DFFQXL \temp78_reg[7]  ( .D(N103), .CK(clk), .Q(temp78[7]) );
  DFFQXL \temp78_reg[6]  ( .D(N102), .CK(clk), .Q(temp78[6]) );
  DFFQXL \temp78_reg[5]  ( .D(N101), .CK(clk), .Q(temp78[5]) );
  DFFQXL \temp1234_reg[13]  ( .D(N141), .CK(clk), .Q(temp1234[13]) );
  DFFQXL \temp1234_reg[12]  ( .D(N140), .CK(clk), .Q(temp1234[12]) );
  DFFQXL \temp1234_reg[11]  ( .D(N139), .CK(clk), .Q(temp1234[11]) );
  DFFQXL \temp1234_reg[10]  ( .D(N138), .CK(clk), .Q(temp1234[10]) );
  DFFQXL \temp1234_reg[9]  ( .D(N137), .CK(clk), .Q(temp1234[9]) );
  DFFQXL \temp1234_reg[8]  ( .D(N136), .CK(clk), .Q(temp1234[8]) );
  DFFQXL \temp1234_reg[7]  ( .D(N135), .CK(clk), .Q(temp1234[7]) );
  DFFQXL \temp1234_reg[6]  ( .D(N134), .CK(clk), .Q(temp1234[6]) );
  DFFQXL \temp9_2_reg[6]  ( .D(temp9[6]), .CK(clk), .Q(temp9_2[6]) );
  DFFQXL \temp9_2_reg[5]  ( .D(temp9[5]), .CK(clk), .Q(temp9_2[5]) );
  DFFQXL \temp9_2_reg[4]  ( .D(temp9[4]), .CK(clk), .Q(temp9_2[4]) );
  DFFQXL \temp9_2_reg[3]  ( .D(temp9[3]), .CK(clk), .Q(temp9_2[3]) );
  DFFQXL \temp9_2_reg[2]  ( .D(temp9[2]), .CK(clk), .Q(temp9_2[2]) );
  DFFQXL \temp9_2_reg[1]  ( .D(temp9[1]), .CK(clk), .Q(temp9_2[1]) );
  DFFQXL \temp12_reg[4]  ( .D(N4), .CK(clk), .Q(temp12[4]) );
  DFFQXL \temp12_reg[3]  ( .D(N3), .CK(clk), .Q(temp12[3]) );
  DFFQXL \temp12_reg[2]  ( .D(N2), .CK(clk), .Q(temp12[2]) );
  DFFQXL \temp12_reg[1]  ( .D(N1), .CK(clk), .Q(temp12[1]) );
  DFFQXL \temp56_reg[4]  ( .D(N68), .CK(clk), .Q(temp56[4]) );
  DFFQXL \temp56_reg[3]  ( .D(N67), .CK(clk), .Q(temp56[3]) );
  DFFQXL \temp56_reg[2]  ( .D(N66), .CK(clk), .Q(temp56[2]) );
  DFFQXL \temp56_reg[1]  ( .D(N65), .CK(clk), .Q(temp56[1]) );
  DFFQXL \temp5678_reg[4]  ( .D(N164), .CK(clk), .Q(temp5678[4]) );
  DFFQXL \temp5678_reg[3]  ( .D(N163), .CK(clk), .Q(temp5678[3]) );
  DFFQXL \temp5678_reg[2]  ( .D(N162), .CK(clk), .Q(temp5678[2]) );
  DFFQXL \temp5678_reg[1]  ( .D(N161), .CK(clk), .Q(temp5678[1]) );
  DFFQXL \temp34_reg[4]  ( .D(N36), .CK(clk), .Q(temp34[4]) );
  DFFQXL \temp34_reg[3]  ( .D(N35), .CK(clk), .Q(temp34[3]) );
  DFFQXL \temp34_reg[2]  ( .D(N34), .CK(clk), .Q(temp34[2]) );
  DFFQXL \temp34_reg[1]  ( .D(N33), .CK(clk), .Q(temp34[1]) );
  DFFQXL \temp78_reg[4]  ( .D(N100), .CK(clk), .Q(temp78[4]) );
  DFFQXL \temp78_reg[3]  ( .D(N99), .CK(clk), .Q(temp78[3]) );
  DFFQXL \temp78_reg[2]  ( .D(N98), .CK(clk), .Q(temp78[2]) );
  DFFQXL \temp78_reg[1]  ( .D(N97), .CK(clk), .Q(temp78[1]) );
  DFFQXL \temp1234_reg[5]  ( .D(N133), .CK(clk), .Q(temp1234[5]) );
  DFFQXL \temp1234_reg[4]  ( .D(N132), .CK(clk), .Q(temp1234[4]) );
  DFFQXL \temp1234_reg[3]  ( .D(N131), .CK(clk), .Q(temp1234[3]) );
  DFFQXL \temp1234_reg[2]  ( .D(N130), .CK(clk), .Q(temp1234[2]) );
  DFFQXL \temp1234_reg[1]  ( .D(N129), .CK(clk), .Q(temp1234[1]) );
  DFFQXL \total_reg[31]  ( .D(N255), .CK(clk), .Q(total[31]) );
  DFFQXL \total_reg[30]  ( .D(N254), .CK(clk), .Q(total[30]) );
  DFFQXL \total_reg[29]  ( .D(N253), .CK(clk), .Q(total[29]) );
  DFFQXL \total_reg[28]  ( .D(N252), .CK(clk), .Q(total[28]) );
  DFFQXL \total_reg[27]  ( .D(N251), .CK(clk), .Q(total[27]) );
  DFFQXL \total_reg[26]  ( .D(N250), .CK(clk), .Q(total[26]) );
  DFFQXL \total_reg[25]  ( .D(N249), .CK(clk), .Q(total[25]) );
  DFFQXL \total_reg[24]  ( .D(N248), .CK(clk), .Q(total[24]) );
  DFFQXL \total_reg[23]  ( .D(N247), .CK(clk), .Q(total[23]) );
  DFFQXL \total_reg[22]  ( .D(N246), .CK(clk), .Q(total[22]) );
  DFFQXL \total_reg[21]  ( .D(N245), .CK(clk), .Q(total[21]) );
  DFFQXL \total_reg[20]  ( .D(N244), .CK(clk), .Q(total[20]) );
  DFFQXL \total_reg[19]  ( .D(N243), .CK(clk), .Q(total[19]) );
  DFFQXL \total_reg[18]  ( .D(N242), .CK(clk), .Q(total[18]) );
  DFFQXL \total_reg[17]  ( .D(N241), .CK(clk), .Q(total[17]) );
  DFFQXL \total_reg[16]  ( .D(N240), .CK(clk), .Q(total[16]) );
  DFFQXL \total_reg[15]  ( .D(N239), .CK(clk), .Q(total[15]) );
  DFFQXL \total_reg[14]  ( .D(N238), .CK(clk), .Q(total[14]) );
  DFFQXL \total_reg[13]  ( .D(N237), .CK(clk), .Q(total[13]) );
  DFFQXL \total_reg[12]  ( .D(N236), .CK(clk), .Q(total[12]) );
  DFFQXL \total_reg[11]  ( .D(N235), .CK(clk), .Q(total[11]) );
  DFFQXL \total_reg[10]  ( .D(N234), .CK(clk), .Q(total[10]) );
  DFFQXL \total_reg[9]  ( .D(N233), .CK(clk), .Q(total[9]) );
  DFFQXL \total_reg[8]  ( .D(N232), .CK(clk), .Q(total[8]) );
  DFFQXL \total_reg[7]  ( .D(N231), .CK(clk), .Q(total[7]) );
  DFFQXL \total_reg[6]  ( .D(N230), .CK(clk), .Q(total[6]) );
  DFFQXL \total_reg[5]  ( .D(N229), .CK(clk), .Q(total[5]) );
  DFFQXL \total_reg[4]  ( .D(N228), .CK(clk), .Q(total[4]) );
  DFFQXL \total_reg[3]  ( .D(N227), .CK(clk), .Q(total[3]) );
  DFFQXL \total_reg[2]  ( .D(N226), .CK(clk), .Q(total[2]) );
  DFFQXL \total_reg[1]  ( .D(N225), .CK(clk), .Q(total[1]) );
  DFFQXL \total_reg[0]  ( .D(N224), .CK(clk), .Q(total[0]) );
  DFFQXL \temp34_reg[0]  ( .D(N32), .CK(clk), .Q(temp34[0]) );
  DFFQXL \temp78_reg[0]  ( .D(N96), .CK(clk), .Q(temp78[0]) );
  DFFQXL \temp1234_reg[0]  ( .D(N128), .CK(clk), .Q(temp1234[0]) );
  DFFQXL \temp12_reg[0]  ( .D(N0), .CK(clk), .Q(temp12[0]) );
  DFFQXL \temp56_reg[0]  ( .D(N64), .CK(clk), .Q(temp56[0]) );
  DFFQXL \temp5678_reg[0]  ( .D(N160), .CK(clk), .Q(temp5678[0]) );
  DFFQXL \temp9_2_reg[0]  ( .D(temp9[0]), .CK(clk), .Q(temp9_2[0]) );
  DFFQXL \temp9_reg[31]  ( .D(in9[31]), .CK(clk), .Q(temp9[31]) );
  DFFQXL \temp9_reg[30]  ( .D(in9[30]), .CK(clk), .Q(temp9[30]) );
  DFFQXL \temp9_reg[29]  ( .D(in9[29]), .CK(clk), .Q(temp9[29]) );
  DFFQXL \temp9_reg[28]  ( .D(in9[28]), .CK(clk), .Q(temp9[28]) );
  DFFQXL \temp9_reg[27]  ( .D(in9[27]), .CK(clk), .Q(temp9[27]) );
  DFFQXL \temp9_reg[26]  ( .D(in9[26]), .CK(clk), .Q(temp9[26]) );
  DFFQXL \temp9_reg[25]  ( .D(in9[25]), .CK(clk), .Q(temp9[25]) );
  DFFQXL \temp9_reg[24]  ( .D(in9[24]), .CK(clk), .Q(temp9[24]) );
  DFFQXL \temp9_reg[23]  ( .D(in9[23]), .CK(clk), .Q(temp9[23]) );
  DFFQXL \temp9_reg[22]  ( .D(in9[22]), .CK(clk), .Q(temp9[22]) );
  DFFQXL \temp9_reg[21]  ( .D(in9[21]), .CK(clk), .Q(temp9[21]) );
  DFFQXL \temp9_reg[20]  ( .D(in9[20]), .CK(clk), .Q(temp9[20]) );
  DFFQXL \temp9_reg[19]  ( .D(in9[19]), .CK(clk), .Q(temp9[19]) );
  DFFQXL \temp9_reg[18]  ( .D(in9[18]), .CK(clk), .Q(temp9[18]) );
  DFFQXL \temp9_reg[17]  ( .D(in9[17]), .CK(clk), .Q(temp9[17]) );
  DFFQXL \temp9_reg[16]  ( .D(in9[16]), .CK(clk), .Q(temp9[16]) );
  DFFQXL \temp9_reg[15]  ( .D(in9[15]), .CK(clk), .Q(temp9[15]) );
  DFFQXL \temp9_reg[14]  ( .D(in9[14]), .CK(clk), .Q(temp9[14]) );
  DFFQXL \temp9_reg[13]  ( .D(in9[13]), .CK(clk), .Q(temp9[13]) );
  DFFQXL \temp9_reg[12]  ( .D(in9[12]), .CK(clk), .Q(temp9[12]) );
  DFFQXL \temp9_reg[11]  ( .D(in9[11]), .CK(clk), .Q(temp9[11]) );
  DFFQXL \temp9_reg[10]  ( .D(in9[10]), .CK(clk), .Q(temp9[10]) );
  DFFQXL \temp9_reg[9]  ( .D(in9[9]), .CK(clk), .Q(temp9[9]) );
  DFFQXL \temp9_reg[8]  ( .D(in9[8]), .CK(clk), .Q(temp9[8]) );
  DFFQXL \temp9_reg[7]  ( .D(in9[7]), .CK(clk), .Q(temp9[7]) );
  DFFQXL \temp9_reg[6]  ( .D(in9[6]), .CK(clk), .Q(temp9[6]) );
  DFFQXL \temp9_reg[5]  ( .D(in9[5]), .CK(clk), .Q(temp9[5]) );
  DFFQXL \temp9_reg[4]  ( .D(in9[4]), .CK(clk), .Q(temp9[4]) );
  DFFQXL \temp9_reg[3]  ( .D(in9[3]), .CK(clk), .Q(temp9[3]) );
  DFFQXL \temp9_reg[2]  ( .D(in9[2]), .CK(clk), .Q(temp9[2]) );
  DFFQXL \temp9_reg[1]  ( .D(in9[1]), .CK(clk), .Q(temp9[1]) );
  DFFQXL \temp9_reg[0]  ( .D(in9[0]), .CK(clk), .Q(temp9[0]) );
endmodule


module Adder_tree_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_tree_1 ( in1, in2, in3, in4, in5, in6, in7, in8, in9, total, clk
 );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  input [31:0] in5;
  input [31:0] in6;
  input [31:0] in7;
  input [31:0] in8;
  input [31:0] in9;
  output [31:0] total;
  input clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N223, N222, N221, N220, N219, N218, N217, N216,
         N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205,
         N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194,
         N193, N192;
  wire   [31:0] temp9;
  wire   [31:0] temp12;
  wire   [31:0] temp34;
  wire   [31:0] temp56;
  wire   [31:0] temp78;
  wire   [31:0] temp1234;
  wire   [31:0] temp5678;
  wire   [31:0] temp9_2;

  Adder_tree_1_DW01_add_0 add_29 ( .A(temp56), .B(temp78), .CI(1'b0), .SUM({
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160}) );
  Adder_tree_1_DW01_add_1 add_28 ( .A(temp12), .B(temp34), .CI(1'b0), .SUM({
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, 
        N135, N134, N133, N132, N131, N130, N129, N128}) );
  Adder_tree_1_DW01_add_2 add_25 ( .A(in7), .B(in8), .CI(1'b0), .SUM({N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96}) );
  Adder_tree_1_DW01_add_3 add_24 ( .A(in5), .B(in6), .CI(1'b0), .SUM({N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64}) );
  Adder_tree_1_DW01_add_4 add_23 ( .A(in3), .B(in4), .CI(1'b0), .SUM({N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32}) );
  Adder_tree_1_DW01_add_5 add_22 ( .A(in1), .B(in2), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Adder_tree_1_DW01_add_7 add_1_root_add_0_root_add_32_2 ( .A(temp9_2), .B(
        temp1234), .CI(1'b0), .SUM({N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 
        N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, 
        N192}) );
  Adder_tree_1_DW01_add_6 add_0_root_add_0_root_add_32_2 ( .A(temp5678), .B({
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192}), .CI(1'b0), .SUM({
        N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, 
        N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, 
        N231, N230, N229, N228, N227, N226, N225, N224}) );
  DFFQXL \temp9_2_reg[31]  ( .D(temp9[31]), .CK(clk), .Q(temp9_2[31]) );
  DFFQXL \temp9_2_reg[30]  ( .D(temp9[30]), .CK(clk), .Q(temp9_2[30]) );
  DFFQXL \temp9_2_reg[29]  ( .D(temp9[29]), .CK(clk), .Q(temp9_2[29]) );
  DFFQXL \temp12_reg[31]  ( .D(N31), .CK(clk), .Q(temp12[31]) );
  DFFQXL \temp12_reg[30]  ( .D(N30), .CK(clk), .Q(temp12[30]) );
  DFFQXL \temp12_reg[29]  ( .D(N29), .CK(clk), .Q(temp12[29]) );
  DFFQXL \temp12_reg[28]  ( .D(N28), .CK(clk), .Q(temp12[28]) );
  DFFQXL \temp12_reg[27]  ( .D(N27), .CK(clk), .Q(temp12[27]) );
  DFFQXL \temp56_reg[31]  ( .D(N95), .CK(clk), .Q(temp56[31]) );
  DFFQXL \temp56_reg[30]  ( .D(N94), .CK(clk), .Q(temp56[30]) );
  DFFQXL \temp56_reg[29]  ( .D(N93), .CK(clk), .Q(temp56[29]) );
  DFFQXL \temp56_reg[28]  ( .D(N92), .CK(clk), .Q(temp56[28]) );
  DFFQXL \temp56_reg[27]  ( .D(N91), .CK(clk), .Q(temp56[27]) );
  DFFQXL \temp5678_reg[31]  ( .D(N191), .CK(clk), .Q(temp5678[31]) );
  DFFQXL \temp5678_reg[30]  ( .D(N190), .CK(clk), .Q(temp5678[30]) );
  DFFQXL \temp5678_reg[29]  ( .D(N189), .CK(clk), .Q(temp5678[29]) );
  DFFQXL \temp5678_reg[28]  ( .D(N188), .CK(clk), .Q(temp5678[28]) );
  DFFQXL \temp5678_reg[27]  ( .D(N187), .CK(clk), .Q(temp5678[27]) );
  DFFQXL \temp34_reg[31]  ( .D(N63), .CK(clk), .Q(temp34[31]) );
  DFFQXL \temp34_reg[30]  ( .D(N62), .CK(clk), .Q(temp34[30]) );
  DFFQXL \temp34_reg[29]  ( .D(N61), .CK(clk), .Q(temp34[29]) );
  DFFQXL \temp34_reg[28]  ( .D(N60), .CK(clk), .Q(temp34[28]) );
  DFFQXL \temp34_reg[27]  ( .D(N59), .CK(clk), .Q(temp34[27]) );
  DFFQXL \temp78_reg[31]  ( .D(N127), .CK(clk), .Q(temp78[31]) );
  DFFQXL \temp78_reg[30]  ( .D(N126), .CK(clk), .Q(temp78[30]) );
  DFFQXL \temp78_reg[29]  ( .D(N125), .CK(clk), .Q(temp78[29]) );
  DFFQXL \temp78_reg[28]  ( .D(N124), .CK(clk), .Q(temp78[28]) );
  DFFQXL \temp78_reg[27]  ( .D(N123), .CK(clk), .Q(temp78[27]) );
  DFFQXL \temp1234_reg[31]  ( .D(N159), .CK(clk), .Q(temp1234[31]) );
  DFFQXL \temp1234_reg[30]  ( .D(N158), .CK(clk), .Q(temp1234[30]) );
  DFFQXL \temp1234_reg[29]  ( .D(N157), .CK(clk), .Q(temp1234[29]) );
  DFFQXL \temp9_2_reg[28]  ( .D(temp9[28]), .CK(clk), .Q(temp9_2[28]) );
  DFFQXL \temp9_2_reg[27]  ( .D(temp9[27]), .CK(clk), .Q(temp9_2[27]) );
  DFFQXL \temp9_2_reg[26]  ( .D(temp9[26]), .CK(clk), .Q(temp9_2[26]) );
  DFFQXL \temp9_2_reg[25]  ( .D(temp9[25]), .CK(clk), .Q(temp9_2[25]) );
  DFFQXL \temp9_2_reg[24]  ( .D(temp9[24]), .CK(clk), .Q(temp9_2[24]) );
  DFFQXL \temp9_2_reg[23]  ( .D(temp9[23]), .CK(clk), .Q(temp9_2[23]) );
  DFFQXL \temp9_2_reg[22]  ( .D(temp9[22]), .CK(clk), .Q(temp9_2[22]) );
  DFFQXL \temp12_reg[26]  ( .D(N26), .CK(clk), .Q(temp12[26]) );
  DFFQXL \temp12_reg[25]  ( .D(N25), .CK(clk), .Q(temp12[25]) );
  DFFQXL \temp12_reg[24]  ( .D(N24), .CK(clk), .Q(temp12[24]) );
  DFFQXL \temp12_reg[23]  ( .D(N23), .CK(clk), .Q(temp12[23]) );
  DFFQXL \temp12_reg[22]  ( .D(N22), .CK(clk), .Q(temp12[22]) );
  DFFQXL \temp12_reg[21]  ( .D(N21), .CK(clk), .Q(temp12[21]) );
  DFFQXL \temp12_reg[20]  ( .D(N20), .CK(clk), .Q(temp12[20]) );
  DFFQXL \temp56_reg[26]  ( .D(N90), .CK(clk), .Q(temp56[26]) );
  DFFQXL \temp56_reg[25]  ( .D(N89), .CK(clk), .Q(temp56[25]) );
  DFFQXL \temp56_reg[24]  ( .D(N88), .CK(clk), .Q(temp56[24]) );
  DFFQXL \temp56_reg[23]  ( .D(N87), .CK(clk), .Q(temp56[23]) );
  DFFQXL \temp56_reg[22]  ( .D(N86), .CK(clk), .Q(temp56[22]) );
  DFFQXL \temp56_reg[21]  ( .D(N85), .CK(clk), .Q(temp56[21]) );
  DFFQXL \temp56_reg[20]  ( .D(N84), .CK(clk), .Q(temp56[20]) );
  DFFQXL \temp5678_reg[26]  ( .D(N186), .CK(clk), .Q(temp5678[26]) );
  DFFQXL \temp5678_reg[25]  ( .D(N185), .CK(clk), .Q(temp5678[25]) );
  DFFQXL \temp5678_reg[24]  ( .D(N184), .CK(clk), .Q(temp5678[24]) );
  DFFQXL \temp5678_reg[23]  ( .D(N183), .CK(clk), .Q(temp5678[23]) );
  DFFQXL \temp5678_reg[22]  ( .D(N182), .CK(clk), .Q(temp5678[22]) );
  DFFQXL \temp5678_reg[21]  ( .D(N181), .CK(clk), .Q(temp5678[21]) );
  DFFQXL \temp5678_reg[20]  ( .D(N180), .CK(clk), .Q(temp5678[20]) );
  DFFQXL \temp34_reg[26]  ( .D(N58), .CK(clk), .Q(temp34[26]) );
  DFFQXL \temp34_reg[25]  ( .D(N57), .CK(clk), .Q(temp34[25]) );
  DFFQXL \temp34_reg[24]  ( .D(N56), .CK(clk), .Q(temp34[24]) );
  DFFQXL \temp34_reg[23]  ( .D(N55), .CK(clk), .Q(temp34[23]) );
  DFFQXL \temp34_reg[22]  ( .D(N54), .CK(clk), .Q(temp34[22]) );
  DFFQXL \temp34_reg[21]  ( .D(N53), .CK(clk), .Q(temp34[21]) );
  DFFQXL \temp34_reg[20]  ( .D(N52), .CK(clk), .Q(temp34[20]) );
  DFFQXL \temp78_reg[26]  ( .D(N122), .CK(clk), .Q(temp78[26]) );
  DFFQXL \temp78_reg[25]  ( .D(N121), .CK(clk), .Q(temp78[25]) );
  DFFQXL \temp78_reg[24]  ( .D(N120), .CK(clk), .Q(temp78[24]) );
  DFFQXL \temp78_reg[23]  ( .D(N119), .CK(clk), .Q(temp78[23]) );
  DFFQXL \temp78_reg[22]  ( .D(N118), .CK(clk), .Q(temp78[22]) );
  DFFQXL \temp78_reg[21]  ( .D(N117), .CK(clk), .Q(temp78[21]) );
  DFFQXL \temp78_reg[20]  ( .D(N116), .CK(clk), .Q(temp78[20]) );
  DFFQXL \temp1234_reg[28]  ( .D(N156), .CK(clk), .Q(temp1234[28]) );
  DFFQXL \temp1234_reg[27]  ( .D(N155), .CK(clk), .Q(temp1234[27]) );
  DFFQXL \temp1234_reg[26]  ( .D(N154), .CK(clk), .Q(temp1234[26]) );
  DFFQXL \temp1234_reg[25]  ( .D(N153), .CK(clk), .Q(temp1234[25]) );
  DFFQXL \temp1234_reg[24]  ( .D(N152), .CK(clk), .Q(temp1234[24]) );
  DFFQXL \temp1234_reg[23]  ( .D(N151), .CK(clk), .Q(temp1234[23]) );
  DFFQXL \temp1234_reg[22]  ( .D(N150), .CK(clk), .Q(temp1234[22]) );
  DFFQXL \temp1234_reg[21]  ( .D(N149), .CK(clk), .Q(temp1234[21]) );
  DFFQXL \temp9_2_reg[21]  ( .D(temp9[21]), .CK(clk), .Q(temp9_2[21]) );
  DFFQXL \temp9_2_reg[20]  ( .D(temp9[20]), .CK(clk), .Q(temp9_2[20]) );
  DFFQXL \temp9_2_reg[19]  ( .D(temp9[19]), .CK(clk), .Q(temp9_2[19]) );
  DFFQXL \temp9_2_reg[18]  ( .D(temp9[18]), .CK(clk), .Q(temp9_2[18]) );
  DFFQXL \temp9_2_reg[17]  ( .D(temp9[17]), .CK(clk), .Q(temp9_2[17]) );
  DFFQXL \temp9_2_reg[16]  ( .D(temp9[16]), .CK(clk), .Q(temp9_2[16]) );
  DFFQXL \temp9_2_reg[15]  ( .D(temp9[15]), .CK(clk), .Q(temp9_2[15]) );
  DFFQXL \temp9_2_reg[14]  ( .D(temp9[14]), .CK(clk), .Q(temp9_2[14]) );
  DFFQXL \temp12_reg[19]  ( .D(N19), .CK(clk), .Q(temp12[19]) );
  DFFQXL \temp12_reg[18]  ( .D(N18), .CK(clk), .Q(temp12[18]) );
  DFFQXL \temp12_reg[17]  ( .D(N17), .CK(clk), .Q(temp12[17]) );
  DFFQXL \temp12_reg[16]  ( .D(N16), .CK(clk), .Q(temp12[16]) );
  DFFQXL \temp12_reg[15]  ( .D(N15), .CK(clk), .Q(temp12[15]) );
  DFFQXL \temp12_reg[14]  ( .D(N14), .CK(clk), .Q(temp12[14]) );
  DFFQXL \temp12_reg[13]  ( .D(N13), .CK(clk), .Q(temp12[13]) );
  DFFQXL \temp12_reg[12]  ( .D(N12), .CK(clk), .Q(temp12[12]) );
  DFFQXL \temp56_reg[19]  ( .D(N83), .CK(clk), .Q(temp56[19]) );
  DFFQXL \temp56_reg[18]  ( .D(N82), .CK(clk), .Q(temp56[18]) );
  DFFQXL \temp56_reg[17]  ( .D(N81), .CK(clk), .Q(temp56[17]) );
  DFFQXL \temp56_reg[16]  ( .D(N80), .CK(clk), .Q(temp56[16]) );
  DFFQXL \temp56_reg[15]  ( .D(N79), .CK(clk), .Q(temp56[15]) );
  DFFQXL \temp56_reg[14]  ( .D(N78), .CK(clk), .Q(temp56[14]) );
  DFFQXL \temp56_reg[13]  ( .D(N77), .CK(clk), .Q(temp56[13]) );
  DFFQXL \temp56_reg[12]  ( .D(N76), .CK(clk), .Q(temp56[12]) );
  DFFQXL \temp5678_reg[19]  ( .D(N179), .CK(clk), .Q(temp5678[19]) );
  DFFQXL \temp5678_reg[18]  ( .D(N178), .CK(clk), .Q(temp5678[18]) );
  DFFQXL \temp5678_reg[17]  ( .D(N177), .CK(clk), .Q(temp5678[17]) );
  DFFQXL \temp5678_reg[16]  ( .D(N176), .CK(clk), .Q(temp5678[16]) );
  DFFQXL \temp5678_reg[15]  ( .D(N175), .CK(clk), .Q(temp5678[15]) );
  DFFQXL \temp5678_reg[14]  ( .D(N174), .CK(clk), .Q(temp5678[14]) );
  DFFQXL \temp5678_reg[13]  ( .D(N173), .CK(clk), .Q(temp5678[13]) );
  DFFQXL \temp5678_reg[12]  ( .D(N172), .CK(clk), .Q(temp5678[12]) );
  DFFQXL \temp34_reg[19]  ( .D(N51), .CK(clk), .Q(temp34[19]) );
  DFFQXL \temp34_reg[18]  ( .D(N50), .CK(clk), .Q(temp34[18]) );
  DFFQXL \temp34_reg[17]  ( .D(N49), .CK(clk), .Q(temp34[17]) );
  DFFQXL \temp34_reg[16]  ( .D(N48), .CK(clk), .Q(temp34[16]) );
  DFFQXL \temp34_reg[15]  ( .D(N47), .CK(clk), .Q(temp34[15]) );
  DFFQXL \temp34_reg[14]  ( .D(N46), .CK(clk), .Q(temp34[14]) );
  DFFQXL \temp34_reg[13]  ( .D(N45), .CK(clk), .Q(temp34[13]) );
  DFFQXL \temp34_reg[12]  ( .D(N44), .CK(clk), .Q(temp34[12]) );
  DFFQXL \temp78_reg[19]  ( .D(N115), .CK(clk), .Q(temp78[19]) );
  DFFQXL \temp78_reg[18]  ( .D(N114), .CK(clk), .Q(temp78[18]) );
  DFFQXL \temp78_reg[17]  ( .D(N113), .CK(clk), .Q(temp78[17]) );
  DFFQXL \temp78_reg[16]  ( .D(N112), .CK(clk), .Q(temp78[16]) );
  DFFQXL \temp78_reg[15]  ( .D(N111), .CK(clk), .Q(temp78[15]) );
  DFFQXL \temp78_reg[14]  ( .D(N110), .CK(clk), .Q(temp78[14]) );
  DFFQXL \temp78_reg[13]  ( .D(N109), .CK(clk), .Q(temp78[13]) );
  DFFQXL \temp78_reg[12]  ( .D(N108), .CK(clk), .Q(temp78[12]) );
  DFFQXL \temp1234_reg[20]  ( .D(N148), .CK(clk), .Q(temp1234[20]) );
  DFFQXL \temp1234_reg[19]  ( .D(N147), .CK(clk), .Q(temp1234[19]) );
  DFFQXL \temp1234_reg[18]  ( .D(N146), .CK(clk), .Q(temp1234[18]) );
  DFFQXL \temp1234_reg[17]  ( .D(N145), .CK(clk), .Q(temp1234[17]) );
  DFFQXL \temp1234_reg[16]  ( .D(N144), .CK(clk), .Q(temp1234[16]) );
  DFFQXL \temp1234_reg[15]  ( .D(N143), .CK(clk), .Q(temp1234[15]) );
  DFFQXL \temp1234_reg[14]  ( .D(N142), .CK(clk), .Q(temp1234[14]) );
  DFFQXL \temp9_2_reg[13]  ( .D(temp9[13]), .CK(clk), .Q(temp9_2[13]) );
  DFFQXL \temp9_2_reg[12]  ( .D(temp9[12]), .CK(clk), .Q(temp9_2[12]) );
  DFFQXL \temp9_2_reg[11]  ( .D(temp9[11]), .CK(clk), .Q(temp9_2[11]) );
  DFFQXL \temp9_2_reg[10]  ( .D(temp9[10]), .CK(clk), .Q(temp9_2[10]) );
  DFFQXL \temp9_2_reg[9]  ( .D(temp9[9]), .CK(clk), .Q(temp9_2[9]) );
  DFFQXL \temp9_2_reg[8]  ( .D(temp9[8]), .CK(clk), .Q(temp9_2[8]) );
  DFFQXL \temp9_2_reg[7]  ( .D(temp9[7]), .CK(clk), .Q(temp9_2[7]) );
  DFFQXL \temp12_reg[11]  ( .D(N11), .CK(clk), .Q(temp12[11]) );
  DFFQXL \temp12_reg[10]  ( .D(N10), .CK(clk), .Q(temp12[10]) );
  DFFQXL \temp12_reg[9]  ( .D(N9), .CK(clk), .Q(temp12[9]) );
  DFFQXL \temp12_reg[8]  ( .D(N8), .CK(clk), .Q(temp12[8]) );
  DFFQXL \temp12_reg[7]  ( .D(N7), .CK(clk), .Q(temp12[7]) );
  DFFQXL \temp12_reg[6]  ( .D(N6), .CK(clk), .Q(temp12[6]) );
  DFFQXL \temp12_reg[5]  ( .D(N5), .CK(clk), .Q(temp12[5]) );
  DFFQXL \temp56_reg[11]  ( .D(N75), .CK(clk), .Q(temp56[11]) );
  DFFQXL \temp56_reg[10]  ( .D(N74), .CK(clk), .Q(temp56[10]) );
  DFFQXL \temp56_reg[9]  ( .D(N73), .CK(clk), .Q(temp56[9]) );
  DFFQXL \temp56_reg[8]  ( .D(N72), .CK(clk), .Q(temp56[8]) );
  DFFQXL \temp56_reg[7]  ( .D(N71), .CK(clk), .Q(temp56[7]) );
  DFFQXL \temp56_reg[6]  ( .D(N70), .CK(clk), .Q(temp56[6]) );
  DFFQXL \temp56_reg[5]  ( .D(N69), .CK(clk), .Q(temp56[5]) );
  DFFQXL \temp5678_reg[11]  ( .D(N171), .CK(clk), .Q(temp5678[11]) );
  DFFQXL \temp5678_reg[10]  ( .D(N170), .CK(clk), .Q(temp5678[10]) );
  DFFQXL \temp5678_reg[9]  ( .D(N169), .CK(clk), .Q(temp5678[9]) );
  DFFQXL \temp5678_reg[8]  ( .D(N168), .CK(clk), .Q(temp5678[8]) );
  DFFQXL \temp5678_reg[7]  ( .D(N167), .CK(clk), .Q(temp5678[7]) );
  DFFQXL \temp5678_reg[6]  ( .D(N166), .CK(clk), .Q(temp5678[6]) );
  DFFQXL \temp5678_reg[5]  ( .D(N165), .CK(clk), .Q(temp5678[5]) );
  DFFQXL \temp34_reg[11]  ( .D(N43), .CK(clk), .Q(temp34[11]) );
  DFFQXL \temp34_reg[10]  ( .D(N42), .CK(clk), .Q(temp34[10]) );
  DFFQXL \temp34_reg[9]  ( .D(N41), .CK(clk), .Q(temp34[9]) );
  DFFQXL \temp34_reg[8]  ( .D(N40), .CK(clk), .Q(temp34[8]) );
  DFFQXL \temp34_reg[7]  ( .D(N39), .CK(clk), .Q(temp34[7]) );
  DFFQXL \temp34_reg[6]  ( .D(N38), .CK(clk), .Q(temp34[6]) );
  DFFQXL \temp34_reg[5]  ( .D(N37), .CK(clk), .Q(temp34[5]) );
  DFFQXL \temp78_reg[11]  ( .D(N107), .CK(clk), .Q(temp78[11]) );
  DFFQXL \temp78_reg[10]  ( .D(N106), .CK(clk), .Q(temp78[10]) );
  DFFQXL \temp78_reg[9]  ( .D(N105), .CK(clk), .Q(temp78[9]) );
  DFFQXL \temp78_reg[8]  ( .D(N104), .CK(clk), .Q(temp78[8]) );
  DFFQXL \temp78_reg[7]  ( .D(N103), .CK(clk), .Q(temp78[7]) );
  DFFQXL \temp78_reg[6]  ( .D(N102), .CK(clk), .Q(temp78[6]) );
  DFFQXL \temp78_reg[5]  ( .D(N101), .CK(clk), .Q(temp78[5]) );
  DFFQXL \temp1234_reg[13]  ( .D(N141), .CK(clk), .Q(temp1234[13]) );
  DFFQXL \temp1234_reg[12]  ( .D(N140), .CK(clk), .Q(temp1234[12]) );
  DFFQXL \temp1234_reg[11]  ( .D(N139), .CK(clk), .Q(temp1234[11]) );
  DFFQXL \temp1234_reg[10]  ( .D(N138), .CK(clk), .Q(temp1234[10]) );
  DFFQXL \temp1234_reg[9]  ( .D(N137), .CK(clk), .Q(temp1234[9]) );
  DFFQXL \temp1234_reg[8]  ( .D(N136), .CK(clk), .Q(temp1234[8]) );
  DFFQXL \temp1234_reg[7]  ( .D(N135), .CK(clk), .Q(temp1234[7]) );
  DFFQXL \temp1234_reg[6]  ( .D(N134), .CK(clk), .Q(temp1234[6]) );
  DFFQXL \temp9_2_reg[6]  ( .D(temp9[6]), .CK(clk), .Q(temp9_2[6]) );
  DFFQXL \temp9_2_reg[5]  ( .D(temp9[5]), .CK(clk), .Q(temp9_2[5]) );
  DFFQXL \temp9_2_reg[4]  ( .D(temp9[4]), .CK(clk), .Q(temp9_2[4]) );
  DFFQXL \temp9_2_reg[3]  ( .D(temp9[3]), .CK(clk), .Q(temp9_2[3]) );
  DFFQXL \temp9_2_reg[2]  ( .D(temp9[2]), .CK(clk), .Q(temp9_2[2]) );
  DFFQXL \temp9_2_reg[1]  ( .D(temp9[1]), .CK(clk), .Q(temp9_2[1]) );
  DFFQXL \temp12_reg[4]  ( .D(N4), .CK(clk), .Q(temp12[4]) );
  DFFQXL \temp12_reg[3]  ( .D(N3), .CK(clk), .Q(temp12[3]) );
  DFFQXL \temp12_reg[2]  ( .D(N2), .CK(clk), .Q(temp12[2]) );
  DFFQXL \temp12_reg[1]  ( .D(N1), .CK(clk), .Q(temp12[1]) );
  DFFQXL \temp56_reg[4]  ( .D(N68), .CK(clk), .Q(temp56[4]) );
  DFFQXL \temp56_reg[3]  ( .D(N67), .CK(clk), .Q(temp56[3]) );
  DFFQXL \temp56_reg[2]  ( .D(N66), .CK(clk), .Q(temp56[2]) );
  DFFQXL \temp56_reg[1]  ( .D(N65), .CK(clk), .Q(temp56[1]) );
  DFFQXL \temp5678_reg[4]  ( .D(N164), .CK(clk), .Q(temp5678[4]) );
  DFFQXL \temp5678_reg[3]  ( .D(N163), .CK(clk), .Q(temp5678[3]) );
  DFFQXL \temp5678_reg[2]  ( .D(N162), .CK(clk), .Q(temp5678[2]) );
  DFFQXL \temp5678_reg[1]  ( .D(N161), .CK(clk), .Q(temp5678[1]) );
  DFFQXL \temp34_reg[4]  ( .D(N36), .CK(clk), .Q(temp34[4]) );
  DFFQXL \temp34_reg[3]  ( .D(N35), .CK(clk), .Q(temp34[3]) );
  DFFQXL \temp34_reg[2]  ( .D(N34), .CK(clk), .Q(temp34[2]) );
  DFFQXL \temp34_reg[1]  ( .D(N33), .CK(clk), .Q(temp34[1]) );
  DFFQXL \temp78_reg[4]  ( .D(N100), .CK(clk), .Q(temp78[4]) );
  DFFQXL \temp78_reg[3]  ( .D(N99), .CK(clk), .Q(temp78[3]) );
  DFFQXL \temp78_reg[2]  ( .D(N98), .CK(clk), .Q(temp78[2]) );
  DFFQXL \temp78_reg[1]  ( .D(N97), .CK(clk), .Q(temp78[1]) );
  DFFQXL \temp1234_reg[5]  ( .D(N133), .CK(clk), .Q(temp1234[5]) );
  DFFQXL \temp1234_reg[4]  ( .D(N132), .CK(clk), .Q(temp1234[4]) );
  DFFQXL \temp1234_reg[3]  ( .D(N131), .CK(clk), .Q(temp1234[3]) );
  DFFQXL \temp1234_reg[2]  ( .D(N130), .CK(clk), .Q(temp1234[2]) );
  DFFQXL \temp1234_reg[1]  ( .D(N129), .CK(clk), .Q(temp1234[1]) );
  DFFQXL \total_reg[31]  ( .D(N255), .CK(clk), .Q(total[31]) );
  DFFQXL \total_reg[30]  ( .D(N254), .CK(clk), .Q(total[30]) );
  DFFQXL \total_reg[29]  ( .D(N253), .CK(clk), .Q(total[29]) );
  DFFQXL \total_reg[28]  ( .D(N252), .CK(clk), .Q(total[28]) );
  DFFQXL \total_reg[27]  ( .D(N251), .CK(clk), .Q(total[27]) );
  DFFQXL \total_reg[26]  ( .D(N250), .CK(clk), .Q(total[26]) );
  DFFQXL \total_reg[25]  ( .D(N249), .CK(clk), .Q(total[25]) );
  DFFQXL \total_reg[24]  ( .D(N248), .CK(clk), .Q(total[24]) );
  DFFQXL \total_reg[23]  ( .D(N247), .CK(clk), .Q(total[23]) );
  DFFQXL \total_reg[22]  ( .D(N246), .CK(clk), .Q(total[22]) );
  DFFQXL \total_reg[21]  ( .D(N245), .CK(clk), .Q(total[21]) );
  DFFQXL \total_reg[20]  ( .D(N244), .CK(clk), .Q(total[20]) );
  DFFQXL \total_reg[19]  ( .D(N243), .CK(clk), .Q(total[19]) );
  DFFQXL \total_reg[18]  ( .D(N242), .CK(clk), .Q(total[18]) );
  DFFQXL \total_reg[17]  ( .D(N241), .CK(clk), .Q(total[17]) );
  DFFQXL \total_reg[16]  ( .D(N240), .CK(clk), .Q(total[16]) );
  DFFQXL \total_reg[15]  ( .D(N239), .CK(clk), .Q(total[15]) );
  DFFQXL \total_reg[14]  ( .D(N238), .CK(clk), .Q(total[14]) );
  DFFQXL \total_reg[13]  ( .D(N237), .CK(clk), .Q(total[13]) );
  DFFQXL \total_reg[12]  ( .D(N236), .CK(clk), .Q(total[12]) );
  DFFQXL \total_reg[11]  ( .D(N235), .CK(clk), .Q(total[11]) );
  DFFQXL \total_reg[10]  ( .D(N234), .CK(clk), .Q(total[10]) );
  DFFQXL \total_reg[9]  ( .D(N233), .CK(clk), .Q(total[9]) );
  DFFQXL \total_reg[8]  ( .D(N232), .CK(clk), .Q(total[8]) );
  DFFQXL \total_reg[7]  ( .D(N231), .CK(clk), .Q(total[7]) );
  DFFQXL \total_reg[6]  ( .D(N230), .CK(clk), .Q(total[6]) );
  DFFQXL \total_reg[5]  ( .D(N229), .CK(clk), .Q(total[5]) );
  DFFQXL \total_reg[4]  ( .D(N228), .CK(clk), .Q(total[4]) );
  DFFQXL \total_reg[3]  ( .D(N227), .CK(clk), .Q(total[3]) );
  DFFQXL \total_reg[2]  ( .D(N226), .CK(clk), .Q(total[2]) );
  DFFQXL \total_reg[1]  ( .D(N225), .CK(clk), .Q(total[1]) );
  DFFQXL \total_reg[0]  ( .D(N224), .CK(clk), .Q(total[0]) );
  DFFQXL \temp34_reg[0]  ( .D(N32), .CK(clk), .Q(temp34[0]) );
  DFFQXL \temp78_reg[0]  ( .D(N96), .CK(clk), .Q(temp78[0]) );
  DFFQXL \temp1234_reg[0]  ( .D(N128), .CK(clk), .Q(temp1234[0]) );
  DFFQXL \temp12_reg[0]  ( .D(N0), .CK(clk), .Q(temp12[0]) );
  DFFQXL \temp56_reg[0]  ( .D(N64), .CK(clk), .Q(temp56[0]) );
  DFFQXL \temp5678_reg[0]  ( .D(N160), .CK(clk), .Q(temp5678[0]) );
  DFFQXL \temp9_2_reg[0]  ( .D(temp9[0]), .CK(clk), .Q(temp9_2[0]) );
  DFFQXL \temp9_reg[31]  ( .D(in9[31]), .CK(clk), .Q(temp9[31]) );
  DFFQXL \temp9_reg[30]  ( .D(in9[30]), .CK(clk), .Q(temp9[30]) );
  DFFQXL \temp9_reg[29]  ( .D(in9[29]), .CK(clk), .Q(temp9[29]) );
  DFFQXL \temp9_reg[28]  ( .D(in9[28]), .CK(clk), .Q(temp9[28]) );
  DFFQXL \temp9_reg[27]  ( .D(in9[27]), .CK(clk), .Q(temp9[27]) );
  DFFQXL \temp9_reg[26]  ( .D(in9[26]), .CK(clk), .Q(temp9[26]) );
  DFFQXL \temp9_reg[25]  ( .D(in9[25]), .CK(clk), .Q(temp9[25]) );
  DFFQXL \temp9_reg[24]  ( .D(in9[24]), .CK(clk), .Q(temp9[24]) );
  DFFQXL \temp9_reg[23]  ( .D(in9[23]), .CK(clk), .Q(temp9[23]) );
  DFFQXL \temp9_reg[22]  ( .D(in9[22]), .CK(clk), .Q(temp9[22]) );
  DFFQXL \temp9_reg[21]  ( .D(in9[21]), .CK(clk), .Q(temp9[21]) );
  DFFQXL \temp9_reg[20]  ( .D(in9[20]), .CK(clk), .Q(temp9[20]) );
  DFFQXL \temp9_reg[19]  ( .D(in9[19]), .CK(clk), .Q(temp9[19]) );
  DFFQXL \temp9_reg[18]  ( .D(in9[18]), .CK(clk), .Q(temp9[18]) );
  DFFQXL \temp9_reg[17]  ( .D(in9[17]), .CK(clk), .Q(temp9[17]) );
  DFFQXL \temp9_reg[16]  ( .D(in9[16]), .CK(clk), .Q(temp9[16]) );
  DFFQXL \temp9_reg[15]  ( .D(in9[15]), .CK(clk), .Q(temp9[15]) );
  DFFQXL \temp9_reg[14]  ( .D(in9[14]), .CK(clk), .Q(temp9[14]) );
  DFFQXL \temp9_reg[13]  ( .D(in9[13]), .CK(clk), .Q(temp9[13]) );
  DFFQXL \temp9_reg[12]  ( .D(in9[12]), .CK(clk), .Q(temp9[12]) );
  DFFQXL \temp9_reg[11]  ( .D(in9[11]), .CK(clk), .Q(temp9[11]) );
  DFFQXL \temp9_reg[10]  ( .D(in9[10]), .CK(clk), .Q(temp9[10]) );
  DFFQXL \temp9_reg[9]  ( .D(in9[9]), .CK(clk), .Q(temp9[9]) );
  DFFQXL \temp9_reg[8]  ( .D(in9[8]), .CK(clk), .Q(temp9[8]) );
  DFFQXL \temp9_reg[7]  ( .D(in9[7]), .CK(clk), .Q(temp9[7]) );
  DFFQXL \temp9_reg[6]  ( .D(in9[6]), .CK(clk), .Q(temp9[6]) );
  DFFQXL \temp9_reg[5]  ( .D(in9[5]), .CK(clk), .Q(temp9[5]) );
  DFFQXL \temp9_reg[4]  ( .D(in9[4]), .CK(clk), .Q(temp9[4]) );
  DFFQXL \temp9_reg[3]  ( .D(in9[3]), .CK(clk), .Q(temp9[3]) );
  DFFQXL \temp9_reg[2]  ( .D(in9[2]), .CK(clk), .Q(temp9[2]) );
  DFFQXL \temp9_reg[1]  ( .D(in9[1]), .CK(clk), .Q(temp9[1]) );
  DFFQXL \temp9_reg[0]  ( .D(in9[0]), .CK(clk), .Q(temp9[0]) );
endmodule


module TOP ( clk, in_pixel, kernal1_00, kernal1_01, kernal1_02, kernal1_10, 
        kernal1_11, kernal1_12, kernal1_20, kernal1_21, kernal1_22, kernal2_00, 
        kernal2_01, kernal2_02, kernal2_10, kernal2_11, kernal2_12, kernal2_20, 
        kernal2_21, kernal2_22, kernal3_00, kernal3_01, kernal3_02, kernal3_10, 
        kernal3_11, kernal3_12, kernal3_20, kernal3_21, kernal3_22, kernal4_00, 
        kernal4_01, kernal4_02, kernal4_10, kernal4_11, kernal4_12, kernal4_20, 
        kernal4_21, kernal4_22, bias1, bias2, bias3, bias4, partial_sum1, 
        partial_sum2, partial_sum3, partial_sum4 );
  input [7:0] in_pixel;
  input [15:0] kernal1_00;
  input [15:0] kernal1_01;
  input [15:0] kernal1_02;
  input [15:0] kernal1_10;
  input [15:0] kernal1_11;
  input [15:0] kernal1_12;
  input [15:0] kernal1_20;
  input [15:0] kernal1_21;
  input [15:0] kernal1_22;
  input [15:0] kernal2_00;
  input [15:0] kernal2_01;
  input [15:0] kernal2_02;
  input [15:0] kernal2_10;
  input [15:0] kernal2_11;
  input [15:0] kernal2_12;
  input [15:0] kernal2_20;
  input [15:0] kernal2_21;
  input [15:0] kernal2_22;
  input [15:0] kernal3_00;
  input [15:0] kernal3_01;
  input [15:0] kernal3_02;
  input [15:0] kernal3_10;
  input [15:0] kernal3_11;
  input [15:0] kernal3_12;
  input [15:0] kernal3_20;
  input [15:0] kernal3_21;
  input [15:0] kernal3_22;
  input [15:0] kernal4_00;
  input [15:0] kernal4_01;
  input [15:0] kernal4_02;
  input [15:0] kernal4_10;
  input [15:0] kernal4_11;
  input [15:0] kernal4_12;
  input [15:0] kernal4_20;
  input [15:0] kernal4_21;
  input [15:0] kernal4_22;
  input [15:0] bias1;
  input [15:0] bias2;
  input [15:0] bias3;
  input [15:0] bias4;
  output [31:0] partial_sum1;
  output [31:0] partial_sum2;
  output [31:0] partial_sum3;
  output [31:0] partial_sum4;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [7:0] pixel_00;
  wire   [7:0] pixel_01;
  wire   [7:0] pixel_02;
  wire   [7:0] pixel_10;
  wire   [7:0] pixel_11;
  wire   [7:0] pixel_12;
  wire   [7:0] pixel_20;
  wire   [7:0] pixel_21;
  wire   [7:0] pixel_22;
  wire   [31:0] out_pixel_pe1;
  wire   [31:0] out_pixel_pe2;
  wire   [31:0] out_pixel_pe3;
  wire   [31:0] out_pixel_pe4;
  wire   [31:0] out_pixel_pe5;
  wire   [31:0] out_pixel_pe6;
  wire   [31:0] out_pixel_pe7;
  wire   [31:0] out_pixel_pe8;
  wire   [31:0] out_pixel_pe9;
  wire   [31:0] out2_pixel_pe1;
  wire   [31:0] out2_pixel_pe2;
  wire   [31:0] out2_pixel_pe3;
  wire   [31:0] out2_pixel_pe4;
  wire   [31:0] out2_pixel_pe5;
  wire   [31:0] out2_pixel_pe6;
  wire   [31:0] out2_pixel_pe7;
  wire   [31:0] out2_pixel_pe8;
  wire   [31:0] out2_pixel_pe9;
  wire   [31:0] out3_pixel_pe1;
  wire   [31:0] out3_pixel_pe2;
  wire   [31:0] out3_pixel_pe3;
  wire   [31:0] out3_pixel_pe4;
  wire   [31:0] out3_pixel_pe5;
  wire   [31:0] out3_pixel_pe6;
  wire   [31:0] out3_pixel_pe7;
  wire   [31:0] out3_pixel_pe8;
  wire   [31:0] out3_pixel_pe9;
  wire   [31:0] out4_pixel_pe1;
  wire   [31:0] out4_pixel_pe2;
  wire   [31:0] out4_pixel_pe3;
  wire   [31:0] out4_pixel_pe4;
  wire   [31:0] out4_pixel_pe5;
  wire   [31:0] out4_pixel_pe6;
  wire   [31:0] out4_pixel_pe7;
  wire   [31:0] out4_pixel_pe8;
  wire   [31:0] out4_pixel_pe9;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287;

  line_buffer LB ( .clk(clk), .pixel_00(pixel_00), .pixel_01(pixel_01), 
        .pixel_02(pixel_02), .pixel_10(pixel_10), .pixel_11(pixel_11), 
        .pixel_12(pixel_12), .pixel_20(pixel_20), .pixel_21(pixel_21), 
        .pixel_22(pixel_22), .in_pixel(in_pixel) );
  PE_0 pe1 ( .pixel_00({n17, pixel_00[6:0]}), .pixel_01({n15, pixel_01[6:0]}), 
        .pixel_02({n13, pixel_02[6:0]}), .pixel_10({n11, pixel_10[6:0]}), 
        .pixel_11({n9, pixel_11[6:0]}), .pixel_12({n7, pixel_12[6:0]}), 
        .pixel_20({n5, pixel_20[6:0]}), .pixel_21({n3, pixel_21[6:0]}), 
        .pixel_22({n1, pixel_22[6:0]}), .weight_00(kernal1_00), .weight_01(
        kernal1_01), .weight_02(kernal1_02), .weight_10(kernal1_10), 
        .weight_11(kernal1_11), .weight_12(kernal1_12), .weight_20(kernal1_20), 
        .weight_21(kernal1_21), .weight_22(kernal1_22), .out_pixel_00({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, out_pixel_pe1[23:0]}), .out_pixel_01({SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        out_pixel_pe2[23:0]}), .out_pixel_02({SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, out_pixel_pe3[23:0]}), .out_pixel_10({
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        out_pixel_pe4[23:0]}), .out_pixel_11({SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, out_pixel_pe5[23:0]}), .out_pixel_12({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        out_pixel_pe6[23:0]}), .out_pixel_20({SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, out_pixel_pe7[23:0]}), .out_pixel_21({
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        out_pixel_pe8[23:0]}), .out_pixel_22({SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, out_pixel_pe9[23:0]}), .clk(clk) );
  PE_3 pe2 ( .pixel_00({n17, pixel_00[6:0]}), .pixel_01({n15, pixel_01[6:0]}), 
        .pixel_02({n13, pixel_02[6:0]}), .pixel_10({n11, pixel_10[6:0]}), 
        .pixel_11({n9, pixel_11[6:0]}), .pixel_12({n7, pixel_12[6:0]}), 
        .pixel_20({n5, pixel_20[6:0]}), .pixel_21({n3, pixel_21[6:0]}), 
        .pixel_22({n1, pixel_22[6:0]}), .weight_00(kernal2_00), .weight_01(
        kernal2_01), .weight_02(kernal2_02), .weight_10(kernal2_10), 
        .weight_11(kernal2_11), .weight_12(kernal2_12), .weight_20(kernal2_20), 
        .weight_21(kernal2_21), .weight_22(kernal2_22), .out_pixel_00({
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        out2_pixel_pe1[23:0]}), .out_pixel_01({SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, out2_pixel_pe2[23:0]}), .out_pixel_02({
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        out2_pixel_pe3[23:0]}), .out_pixel_10({SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, out2_pixel_pe4[23:0]}), .out_pixel_11({
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        out2_pixel_pe5[23:0]}), .out_pixel_12({SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, out2_pixel_pe6[23:0]}), .out_pixel_20({
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        out2_pixel_pe7[23:0]}), .out_pixel_21({SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, out2_pixel_pe8[23:0]}), .out_pixel_22({
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        out2_pixel_pe9[23:0]}), .clk(clk) );
  PE_2 pe3 ( .pixel_00({n17, pixel_00[6:0]}), .pixel_01({n15, pixel_01[6:0]}), 
        .pixel_02({n13, pixel_02[6:0]}), .pixel_10({n11, pixel_10[6:0]}), 
        .pixel_11({n9, pixel_11[6:0]}), .pixel_12({n7, pixel_12[6:0]}), 
        .pixel_20({n5, pixel_20[6:0]}), .pixel_21({n3, pixel_21[6:0]}), 
        .pixel_22({n1, pixel_22[6:0]}), .weight_00(kernal3_00), .weight_01(
        kernal3_01), .weight_02(kernal3_02), .weight_10(kernal3_10), 
        .weight_11(kernal3_11), .weight_12(kernal3_12), .weight_20(kernal3_20), 
        .weight_21(kernal3_21), .weight_22(kernal3_22), .out_pixel_00({
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        out3_pixel_pe1[23:0]}), .out_pixel_01({SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, out3_pixel_pe2[23:0]}), .out_pixel_02({
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        out3_pixel_pe3[23:0]}), .out_pixel_10({SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, out3_pixel_pe4[23:0]}), .out_pixel_11({
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        out3_pixel_pe5[23:0]}), .out_pixel_12({SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, 
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, 
        SYNOPSYS_UNCONNECTED__191, out3_pixel_pe6[23:0]}), .out_pixel_20({
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        out3_pixel_pe7[23:0]}), .out_pixel_21({SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, 
        SYNOPSYS_UNCONNECTED__207, out3_pixel_pe8[23:0]}), .out_pixel_22({
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        out3_pixel_pe9[23:0]}), .clk(clk) );
  PE_1 pe4 ( .pixel_00({n17, pixel_00[6:0]}), .pixel_01({n15, pixel_01[6:0]}), 
        .pixel_02({n13, pixel_02[6:0]}), .pixel_10({n11, pixel_10[6:0]}), 
        .pixel_11({n9, pixel_11[6:0]}), .pixel_12({n7, pixel_12[6:0]}), 
        .pixel_20({n5, pixel_20[6:0]}), .pixel_21({n3, pixel_21[6:0]}), 
        .pixel_22({n1, pixel_22[6:0]}), .weight_00(kernal4_00), .weight_01(
        kernal4_01), .weight_02(kernal4_02), .weight_10(kernal4_10), 
        .weight_11(kernal4_11), .weight_12(kernal4_12), .weight_20(kernal4_20), 
        .weight_21(kernal4_21), .weight_22(kernal4_22), .out_pixel_00({
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        out4_pixel_pe1[23:0]}), .out_pixel_01({SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, 
        SYNOPSYS_UNCONNECTED__227, SYNOPSYS_UNCONNECTED__228, 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, out4_pixel_pe2[23:0]}), .out_pixel_02({
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        out4_pixel_pe3[23:0]}), .out_pixel_10({SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, 
        SYNOPSYS_UNCONNECTED__247, out4_pixel_pe4[23:0]}), .out_pixel_11({
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        out4_pixel_pe5[23:0]}), .out_pixel_12({SYNOPSYS_UNCONNECTED__256, 
        SYNOPSYS_UNCONNECTED__257, SYNOPSYS_UNCONNECTED__258, 
        SYNOPSYS_UNCONNECTED__259, SYNOPSYS_UNCONNECTED__260, 
        SYNOPSYS_UNCONNECTED__261, SYNOPSYS_UNCONNECTED__262, 
        SYNOPSYS_UNCONNECTED__263, out4_pixel_pe6[23:0]}), .out_pixel_20({
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        out4_pixel_pe7[23:0]}), .out_pixel_21({SYNOPSYS_UNCONNECTED__272, 
        SYNOPSYS_UNCONNECTED__273, SYNOPSYS_UNCONNECTED__274, 
        SYNOPSYS_UNCONNECTED__275, SYNOPSYS_UNCONNECTED__276, 
        SYNOPSYS_UNCONNECTED__277, SYNOPSYS_UNCONNECTED__278, 
        SYNOPSYS_UNCONNECTED__279, out4_pixel_pe8[23:0]}), .out_pixel_22({
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        out4_pixel_pe9[23:0]}), .clk(clk) );
  Adder_tree_0 adder_tree1 ( .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out_pixel_pe1[23:0]}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, out_pixel_pe2[23:0]}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, out_pixel_pe3[23:0]}), .in4({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, out_pixel_pe4[23:0]}), .in5({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_pixel_pe5[23:0]}), .in6({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_pixel_pe6[23:0]}), .in7({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_pixel_pe7[23:0]}), .in8(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_pixel_pe8[23:0]}), 
        .in9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        out_pixel_pe9[23:0]}), .total(partial_sum1), .clk(clk) );
  Adder_tree_3 adder_tree2 ( .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out2_pixel_pe1[23:0]}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, out2_pixel_pe2[23:0]}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, out2_pixel_pe3[23:0]}), .in4({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, out2_pixel_pe4[23:0]}), .in5({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out2_pixel_pe5[23:0]}), .in6({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out2_pixel_pe6[23:0]}), .in7({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out2_pixel_pe7[23:0]}), 
        .in8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        out2_pixel_pe8[23:0]}), .in9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out2_pixel_pe9[23:0]}), .total(partial_sum2), .clk(clk) );
  Adder_tree_2 adder_tree3 ( .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out3_pixel_pe1[23:0]}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, out3_pixel_pe2[23:0]}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, out3_pixel_pe3[23:0]}), .in4({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, out3_pixel_pe4[23:0]}), .in5({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out3_pixel_pe5[23:0]}), .in6({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out3_pixel_pe6[23:0]}), .in7({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out3_pixel_pe7[23:0]}), 
        .in8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        out3_pixel_pe8[23:0]}), .in9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out3_pixel_pe9[23:0]}), .total(partial_sum3), .clk(clk) );
  Adder_tree_1 adder_tree4 ( .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out4_pixel_pe1[23:0]}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, out4_pixel_pe2[23:0]}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, out4_pixel_pe3[23:0]}), .in4({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, out4_pixel_pe4[23:0]}), .in5({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out4_pixel_pe5[23:0]}), .in6({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out4_pixel_pe6[23:0]}), .in7({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out4_pixel_pe7[23:0]}), 
        .in8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        out4_pixel_pe8[23:0]}), .in9({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out4_pixel_pe9[23:0]}), .total(partial_sum4), .clk(clk) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(pixel_22[7]), .Y(n2) );
  INVX2 U3 ( .A(n4), .Y(n3) );
  INVX2 U4 ( .A(pixel_21[7]), .Y(n4) );
  INVX2 U5 ( .A(n6), .Y(n5) );
  INVX2 U6 ( .A(pixel_20[7]), .Y(n6) );
  INVX2 U7 ( .A(n8), .Y(n7) );
  INVX2 U8 ( .A(pixel_12[7]), .Y(n8) );
  INVX2 U9 ( .A(n10), .Y(n9) );
  INVX2 U10 ( .A(pixel_11[7]), .Y(n10) );
  INVX2 U11 ( .A(n12), .Y(n11) );
  INVX2 U12 ( .A(pixel_10[7]), .Y(n12) );
  INVX2 U13 ( .A(n14), .Y(n13) );
  INVX2 U14 ( .A(pixel_02[7]), .Y(n14) );
  INVX2 U15 ( .A(n16), .Y(n15) );
  INVX2 U16 ( .A(pixel_01[7]), .Y(n16) );
  INVX2 U17 ( .A(n18), .Y(n17) );
  INVX2 U18 ( .A(pixel_00[7]), .Y(n18) );
endmodule

